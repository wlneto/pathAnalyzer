// Benchmark "iscas20_aigs/mem_ctrl" written by ABC on Wed Jan  8 15:30:41 2020

module mem_ctrl  ( clock, 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151  );
  input  clock;
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151;
  reg lo0000, lo0001, lo0002, lo0003, lo0004, lo0005, lo0006, lo0007,
    lo0008, lo0009, lo0010, lo0011, lo0012, lo0013, lo0014, lo0015, lo0016,
    lo0017, lo0018, lo0019, lo0020, lo0021, lo0022, lo0023, lo0024, lo0025,
    lo0026, lo0027, lo0028, lo0029, lo0030, lo0031, lo0032, lo0033, lo0034,
    lo0035, lo0036, lo0037, lo0038, lo0039, lo0040, lo0041, lo0042, lo0043,
    lo0044, lo0045, lo0046, lo0047, lo0048, lo0049, lo0050, lo0051, lo0052,
    lo0053, lo0054, lo0055, lo0056, lo0057, lo0058, lo0059, lo0060, lo0061,
    lo0062, lo0063, lo0064, lo0065, lo0066, lo0067, lo0068, lo0069, lo0070,
    lo0071, lo0072, lo0073, lo0074, lo0075, lo0076, lo0077, lo0078, lo0079,
    lo0080, lo0081, lo0082, lo0083, lo0084, lo0085, lo0086, lo0087, lo0088,
    lo0089, lo0090, lo0091, lo0092, lo0093, lo0094, lo0095, lo0096, lo0097,
    lo0098, lo0099, lo0100, lo0101, lo0102, lo0103, lo0104, lo0105, lo0106,
    lo0107, lo0108, lo0109, lo0110, lo0111, lo0112, lo0113, lo0114, lo0115,
    lo0116, lo0117, lo0118, lo0119, lo0120, lo0121, lo0122, lo0123, lo0124,
    lo0125, lo0126, lo0127, lo0128, lo0129, lo0130, lo0131, lo0132, lo0133,
    lo0134, lo0135, lo0136, lo0137, lo0138, lo0139, lo0140, lo0141, lo0142,
    lo0143, lo0144, lo0145, lo0146, lo0147, lo0148, lo0149, lo0150, lo0151,
    lo0152, lo0153, lo0154, lo0155, lo0156, lo0157, lo0158, lo0159, lo0160,
    lo0161, lo0162, lo0163, lo0164, lo0165, lo0166, lo0167, lo0168, lo0169,
    lo0170, lo0171, lo0172, lo0173, lo0174, lo0175, lo0176, lo0177, lo0178,
    lo0179, lo0180, lo0181, lo0182, lo0183, lo0184, lo0185, lo0186, lo0187,
    lo0188, lo0189, lo0190, lo0191, lo0192, lo0193, lo0194, lo0195, lo0196,
    lo0197, lo0198, lo0199, lo0200, lo0201, lo0202, lo0203, lo0204, lo0205,
    lo0206, lo0207, lo0208, lo0209, lo0210, lo0211, lo0212, lo0213, lo0214,
    lo0215, lo0216, lo0217, lo0218, lo0219, lo0220, lo0221, lo0222, lo0223,
    lo0224, lo0225, lo0226, lo0227, lo0228, lo0229, lo0230, lo0231, lo0232,
    lo0233, lo0234, lo0235, lo0236, lo0237, lo0238, lo0239, lo0240, lo0241,
    lo0242, lo0243, lo0244, lo0245, lo0246, lo0247, lo0248, lo0249, lo0250,
    lo0251, lo0252, lo0253, lo0254, lo0255, lo0256, lo0257, lo0258, lo0259,
    lo0260, lo0261, lo0262, lo0263, lo0264, lo0265, lo0266, lo0267, lo0268,
    lo0269, lo0270, lo0271, lo0272, lo0273, lo0274, lo0275, lo0276, lo0277,
    lo0278, lo0279, lo0280, lo0281, lo0282, lo0283, lo0284, lo0285, lo0286,
    lo0287, lo0288, lo0289, lo0290, lo0291, lo0292, lo0293, lo0294, lo0295,
    lo0296, lo0297, lo0298, lo0299, lo0300, lo0301, lo0302, lo0303, lo0304,
    lo0305, lo0306, lo0307, lo0308, lo0309, lo0310, lo0311, lo0312, lo0313,
    lo0314, lo0315, lo0316, lo0317, lo0318, lo0319, lo0320, lo0321, lo0322,
    lo0323, lo0324, lo0325, lo0326, lo0327, lo0328, lo0329, lo0330, lo0331,
    lo0332, lo0333, lo0334, lo0335, lo0336, lo0337, lo0338, lo0339, lo0340,
    lo0341, lo0342, lo0343, lo0344, lo0345, lo0346, lo0347, lo0348, lo0349,
    lo0350, lo0351, lo0352, lo0353, lo0354, lo0355, lo0356, lo0357, lo0358,
    lo0359, lo0360, lo0361, lo0362, lo0363, lo0364, lo0365, lo0366, lo0367,
    lo0368, lo0369, lo0370, lo0371, lo0372, lo0373, lo0374, lo0375, lo0376,
    lo0377, lo0378, lo0379, lo0380, lo0381, lo0382, lo0383, lo0384, lo0385,
    lo0386, lo0387, lo0388, lo0389, lo0390, lo0391, lo0392, lo0393, lo0394,
    lo0395, lo0396, lo0397, lo0398, lo0399, lo0400, lo0401, lo0402, lo0403,
    lo0404, lo0405, lo0406, lo0407, lo0408, lo0409, lo0410, lo0411, lo0412,
    lo0413, lo0414, lo0415, lo0416, lo0417, lo0418, lo0419, lo0420, lo0421,
    lo0422, lo0423, lo0424, lo0425, lo0426, lo0427, lo0428, lo0429, lo0430,
    lo0431, lo0432, lo0433, lo0434, lo0435, lo0436, lo0437, lo0438, lo0439,
    lo0440, lo0441, lo0442, lo0443, lo0444, lo0445, lo0446, lo0447, lo0448,
    lo0449, lo0450, lo0451, lo0452, lo0453, lo0454, lo0455, lo0456, lo0457,
    lo0458, lo0459, lo0460, lo0461, lo0462, lo0463, lo0464, lo0465, lo0466,
    lo0467, lo0468, lo0469, lo0470, lo0471, lo0472, lo0473, lo0474, lo0475,
    lo0476, lo0477, lo0478, lo0479, lo0480, lo0481, lo0482, lo0483, lo0484,
    lo0485, lo0486, lo0487, lo0488, lo0489, lo0490, lo0491, lo0492, lo0493,
    lo0494, lo0495, lo0496, lo0497, lo0498, lo0499, lo0500, lo0501, lo0502,
    lo0503, lo0504, lo0505, lo0506, lo0507, lo0508, lo0509, lo0510, lo0511,
    lo0512, lo0513, lo0514, lo0515, lo0516, lo0517, lo0518, lo0519, lo0520,
    lo0521, lo0522, lo0523, lo0524, lo0525, lo0526, lo0527, lo0528, lo0529,
    lo0530, lo0531, lo0532, lo0533, lo0534, lo0535, lo0536, lo0537, lo0538,
    lo0539, lo0540, lo0541, lo0542, lo0543, lo0544, lo0545, lo0546, lo0547,
    lo0548, lo0549, lo0550, lo0551, lo0552, lo0553, lo0554, lo0555, lo0556,
    lo0557, lo0558, lo0559, lo0560, lo0561, lo0562, lo0563, lo0564, lo0565,
    lo0566, lo0567, lo0568, lo0569, lo0570, lo0571, lo0572, lo0573, lo0574,
    lo0575, lo0576, lo0577, lo0578, lo0579, lo0580, lo0581, lo0582, lo0583,
    lo0584, lo0585, lo0586, lo0587, lo0588, lo0589, lo0590, lo0591, lo0592,
    lo0593, lo0594, lo0595, lo0596, lo0597, lo0598, lo0599, lo0600, lo0601,
    lo0602, lo0603, lo0604, lo0605, lo0606, lo0607, lo0608, lo0609, lo0610,
    lo0611, lo0612, lo0613, lo0614, lo0615, lo0616, lo0617, lo0618, lo0619,
    lo0620, lo0621, lo0622, lo0623, lo0624, lo0625, lo0626, lo0627, lo0628,
    lo0629, lo0630, lo0631, lo0632, lo0633, lo0634, lo0635, lo0636, lo0637,
    lo0638, lo0639, lo0640, lo0641, lo0642, lo0643, lo0644, lo0645, lo0646,
    lo0647, lo0648, lo0649, lo0650, lo0651, lo0652, lo0653, lo0654, lo0655,
    lo0656, lo0657, lo0658, lo0659, lo0660, lo0661, lo0662, lo0663, lo0664,
    lo0665, lo0666, lo0667, lo0668, lo0669, lo0670, lo0671, lo0672, lo0673,
    lo0674, lo0675, lo0676, lo0677, lo0678, lo0679, lo0680, lo0681, lo0682,
    lo0683, lo0684, lo0685, lo0686, lo0687, lo0688, lo0689, lo0690, lo0691,
    lo0692, lo0693, lo0694, lo0695, lo0696, lo0697, lo0698, lo0699, lo0700,
    lo0701, lo0702, lo0703, lo0704, lo0705, lo0706, lo0707, lo0708, lo0709,
    lo0710, lo0711, lo0712, lo0713, lo0714, lo0715, lo0716, lo0717, lo0718,
    lo0719, lo0720, lo0721, lo0722, lo0723, lo0724, lo0725, lo0726, lo0727,
    lo0728, lo0729, lo0730, lo0731, lo0732, lo0733, lo0734, lo0735, lo0736,
    lo0737, lo0738, lo0739, lo0740, lo0741, lo0742, lo0743, lo0744, lo0745,
    lo0746, lo0747, lo0748, lo0749, lo0750, lo0751, lo0752, lo0753, lo0754,
    lo0755, lo0756, lo0757, lo0758, lo0759, lo0760, lo0761, lo0762, lo0763,
    lo0764, lo0765, lo0766, lo0767, lo0768, lo0769, lo0770, lo0771, lo0772,
    lo0773, lo0774, lo0775, lo0776, lo0777, lo0778, lo0779, lo0780, lo0781,
    lo0782, lo0783, lo0784, lo0785, lo0786, lo0787, lo0788, lo0789, lo0790,
    lo0791, lo0792, lo0793, lo0794, lo0795, lo0796, lo0797, lo0798, lo0799,
    lo0800, lo0801, lo0802, lo0803, lo0804, lo0805, lo0806, lo0807, lo0808,
    lo0809, lo0810, lo0811, lo0812, lo0813, lo0814, lo0815, lo0816, lo0817,
    lo0818, lo0819, lo0820, lo0821, lo0822, lo0823, lo0824, lo0825, lo0826,
    lo0827, lo0828, lo0829, lo0830, lo0831, lo0832, lo0833, lo0834, lo0835,
    lo0836, lo0837, lo0838, lo0839, lo0840, lo0841, lo0842, lo0843, lo0844,
    lo0845, lo0846, lo0847, lo0848, lo0849, lo0850, lo0851, lo0852, lo0853,
    lo0854, lo0855, lo0856, lo0857, lo0858, lo0859, lo0860, lo0861, lo0862,
    lo0863, lo0864, lo0865, lo0866, lo0867, lo0868, lo0869, lo0870, lo0871,
    lo0872, lo0873, lo0874, lo0875, lo0876, lo0877, lo0878, lo0879, lo0880,
    lo0881, lo0882, lo0883, lo0884, lo0885, lo0886, lo0887, lo0888, lo0889,
    lo0890, lo0891, lo0892, lo0893, lo0894, lo0895, lo0896, lo0897, lo0898,
    lo0899, lo0900, lo0901, lo0902, lo0903, lo0904, lo0905, lo0906, lo0907,
    lo0908, lo0909, lo0910, lo0911, lo0912, lo0913, lo0914, lo0915, lo0916,
    lo0917, lo0918, lo0919, lo0920, lo0921, lo0922, lo0923, lo0924, lo0925,
    lo0926, lo0927, lo0928, lo0929, lo0930, lo0931, lo0932, lo0933, lo0934,
    lo0935, lo0936, lo0937, lo0938, lo0939, lo0940, lo0941, lo0942, lo0943,
    lo0944, lo0945, lo0946, lo0947, lo0948, lo0949, lo0950, lo0951, lo0952,
    lo0953, lo0954, lo0955, lo0956, lo0957, lo0958, lo0959, lo0960, lo0961,
    lo0962, lo0963, lo0964, lo0965, lo0966, lo0967, lo0968, lo0969, lo0970,
    lo0971, lo0972, lo0973, lo0974, lo0975, lo0976, lo0977, lo0978, lo0979,
    lo0980, lo0981, lo0982, lo0983, lo0984, lo0985, lo0986, lo0987, lo0988,
    lo0989, lo0990, lo0991, lo0992, lo0993, lo0994, lo0995, lo0996, lo0997,
    lo0998, lo0999, lo1000, lo1001, lo1002, lo1003, lo1004, lo1005, lo1006,
    lo1007, lo1008, lo1009, lo1010, lo1011, lo1012, lo1013, lo1014, lo1015,
    lo1016, lo1017, lo1018, lo1019, lo1020, lo1021, lo1022, lo1023, lo1024,
    lo1025, lo1026, lo1027, lo1028, lo1029, lo1030, lo1031, lo1032, lo1033,
    lo1034, lo1035, lo1036, lo1037, lo1038, lo1039, lo1040, lo1041, lo1042,
    lo1043, lo1044, lo1045, lo1046, lo1047, lo1048, lo1049, lo1050, lo1051,
    lo1052, lo1053, lo1054, lo1055, lo1056, lo1057, lo1058, lo1059, lo1060,
    lo1061, lo1062, lo1063, lo1064, lo1065, lo1066, lo1067, lo1068, lo1069,
    lo1070, lo1071, lo1072, lo1073, lo1074, lo1075, lo1076, lo1077, lo1078,
    lo1079, lo1080, lo1081, lo1082;
  wire new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_,
    new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_,
    new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_,
    new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_,
    new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_,
    new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_,
    new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_,
    new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_,
    new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_,
    new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_,
    new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_,
    new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_,
    new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_,
    new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_,
    new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_,
    new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_,
    new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_,
    new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_,
    new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_,
    new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_,
    new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_,
    new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_,
    new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_,
    new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_,
    new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3666_, new_n3667_,
    new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_,
    new_n3674_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3682_,
    new_n3685_, new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_,
    new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_,
    new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_,
    new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_,
    new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_,
    new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_,
    new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_,
    new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_,
    new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_,
    new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_,
    new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_,
    new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_,
    new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_,
    new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_,
    new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_,
    new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_,
    new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_,
    new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_,
    new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_,
    new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_,
    new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_,
    new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_,
    new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_,
    new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_,
    new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_,
    new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_,
    new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_,
    new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_,
    new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_,
    new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_,
    new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_,
    new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_,
    new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_,
    new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_,
    new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_,
    new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_,
    new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3920_,
    new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_,
    new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_,
    new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_,
    new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_,
    new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_,
    new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_,
    new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_,
    new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_,
    new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_,
    new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_,
    new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_,
    new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_,
    new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_,
    new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_,
    new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_,
    new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_,
    new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_,
    new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_,
    new_n4029_, new_n4030_, new_n4032_, new_n4033_, new_n4034_, new_n4035_,
    new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_,
    new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_,
    new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_,
    new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_,
    new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_,
    new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_,
    new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4148_, new_n4149_, new_n4150_,
    new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_,
    new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_,
    new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_,
    new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_,
    new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_,
    new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_,
    new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_,
    new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_,
    new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_,
    new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_,
    new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_,
    new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_,
    new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_,
    new_n4229_, new_n4230_, new_n4231_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_,
    new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_,
    new_n4274_, new_n4275_, new_n4277_, new_n4278_, new_n4279_, new_n4280_,
    new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_,
    new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_,
    new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4311_, new_n4312_,
    new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_,
    new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_,
    new_n4325_, new_n4326_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_,
    new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_,
    new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4379_, new_n4380_, new_n4381_, new_n4382_,
    new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4388_,
    new_n4389_, new_n4390_, new_n4391_, new_n4393_, new_n4394_, new_n4395_,
    new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_,
    new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4407_, new_n4408_,
    new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_,
    new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4523_, new_n4524_,
    new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_,
    new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_,
    new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_,
    new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_,
    new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_,
    new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_,
    new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_,
    new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_,
    new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_,
    new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_,
    new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_,
    new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4597_,
    new_n4598_, new_n4599_, new_n4602_, new_n4604_, new_n4606_, new_n4608_,
    new_n4610_, new_n4612_, new_n4614_, new_n4615_, new_n4617_, new_n4618_,
    new_n4619_, new_n4620_, new_n4622_, new_n4623_, new_n4625_, new_n4626_,
    new_n4628_, new_n4629_, new_n4631_, new_n4632_, new_n4633_, new_n4634_,
    new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_,
    new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_,
    new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_,
    new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_,
    new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_,
    new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_,
    new_n4671_, new_n4672_, new_n4673_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_,
    new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_,
    new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_,
    new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_,
    new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_,
    new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_,
    new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_,
    new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_,
    new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_,
    new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_,
    new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_,
    new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_,
    new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_,
    new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_,
    new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_,
    new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_,
    new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_,
    new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_,
    new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_,
    new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_,
    new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_,
    new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_,
    new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_,
    new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_,
    new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_,
    new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_,
    new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_,
    new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_,
    new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_,
    new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_,
    new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_,
    new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_,
    new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_,
    new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_,
    new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_,
    new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_,
    new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_,
    new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_,
    new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_,
    new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_,
    new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_,
    new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_,
    new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_,
    new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_,
    new_n5056_, new_n5057_, new_n5058_, new_n5060_, new_n5061_, new_n5062_,
    new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_,
    new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_,
    new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_,
    new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_,
    new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_,
    new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_,
    new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_,
    new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_,
    new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_,
    new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_,
    new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_,
    new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_,
    new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_,
    new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_,
    new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_,
    new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_,
    new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_,
    new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_,
    new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_,
    new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_,
    new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_,
    new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_,
    new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_,
    new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_,
    new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_,
    new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_,
    new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_,
    new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_,
    new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_,
    new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_,
    new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_,
    new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_,
    new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_,
    new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_,
    new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_,
    new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5376_, new_n5377_, new_n5378_,
    new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_,
    new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_,
    new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_,
    new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_,
    new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_,
    new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_,
    new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_,
    new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_,
    new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_,
    new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_,
    new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_,
    new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_,
    new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_,
    new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_,
    new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_,
    new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_,
    new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_,
    new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_,
    new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_,
    new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_,
    new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_,
    new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5511_,
    new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_,
    new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_,
    new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_,
    new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_,
    new_n5536_, new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_,
    new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_,
    new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_,
    new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_,
    new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_,
    new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_,
    new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_,
    new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_,
    new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_,
    new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_,
    new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_,
    new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_,
    new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_,
    new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_,
    new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_,
    new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_,
    new_n5632_, new_n5633_, new_n5634_, new_n5636_, new_n5637_, new_n5638_,
    new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_,
    new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_,
    new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_,
    new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_,
    new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_,
    new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_,
    new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_,
    new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_,
    new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_,
    new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_,
    new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_,
    new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_,
    new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_,
    new_n5717_, new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_,
    new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_,
    new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_,
    new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_,
    new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_,
    new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_,
    new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_,
    new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_,
    new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_,
    new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5898_,
    new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_,
    new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_,
    new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_,
    new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_,
    new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_,
    new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_,
    new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_,
    new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_,
    new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_,
    new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_,
    new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_,
    new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_,
    new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_,
    new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_,
    new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_,
    new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_,
    new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_,
    new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_,
    new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_,
    new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_,
    new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6026_,
    new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_,
    new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_,
    new_n6039_, new_n6040_, new_n6041_, new_n6043_, new_n6044_, new_n6045_,
    new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_,
    new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_,
    new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_, new_n6074_, new_n6075_, new_n6076_,
    new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_,
    new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_,
    new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_,
    new_n6095_, new_n6096_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6106_, new_n6107_, new_n6108_,
    new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_,
    new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_,
    new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_,
    new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_,
    new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_,
    new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_,
    new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_,
    new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_,
    new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_,
    new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_,
    new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_,
    new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_,
    new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_,
    new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_,
    new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_,
    new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_,
    new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_,
    new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_,
    new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_,
    new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_,
    new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_,
    new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_,
    new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_,
    new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_,
    new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_,
    new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_,
    new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_,
    new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_,
    new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_,
    new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_, new_n6289_,
    new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_,
    new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_, new_n6301_,
    new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_, new_n6307_,
    new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_,
    new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_,
    new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_,
    new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_,
    new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_,
    new_n6338_, new_n6340_, new_n6341_, new_n6342_, new_n6343_, new_n6344_,
    new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_, new_n6350_,
    new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_, new_n6356_,
    new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_, new_n6362_,
    new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_, new_n6368_,
    new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_, new_n6374_,
    new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_, new_n6380_,
    new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_, new_n6386_,
    new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_, new_n6392_,
    new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_, new_n6398_,
    new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_, new_n6404_,
    new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_, new_n6410_,
    new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_, new_n6416_,
    new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_, new_n6422_,
    new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_, new_n6428_,
    new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_, new_n6434_,
    new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_, new_n6440_,
    new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_, new_n6446_,
    new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_,
    new_n6453_, new_n6454_, new_n6455_, new_n6457_, new_n6458_, new_n6459_,
    new_n6460_, new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_,
    new_n6466_, new_n6467_, new_n6468_, new_n6469_, new_n6470_, new_n6471_,
    new_n6472_, new_n6473_, new_n6474_, new_n6475_, new_n6476_, new_n6477_,
    new_n6478_, new_n6479_, new_n6480_, new_n6481_, new_n6482_, new_n6483_,
    new_n6484_, new_n6485_, new_n6486_, new_n6487_, new_n6488_, new_n6489_,
    new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_,
    new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_,
    new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_,
    new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_, new_n6513_,
    new_n6514_, new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_,
    new_n6520_, new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_,
    new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_,
    new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_,
    new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_,
    new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_,
    new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_,
    new_n6556_, new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_,
    new_n6562_, new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_,
    new_n6568_, new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_,
    new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_,
    new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_,
    new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_,
    new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_,
    new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_,
    new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_,
    new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_,
    new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_,
    new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_,
    new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_,
    new_n6635_, new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_,
    new_n6641_, new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_,
    new_n6647_, new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_,
    new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_,
    new_n6659_, new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_,
    new_n6665_, new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_,
    new_n6671_, new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_,
    new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_,
    new_n6683_, new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_,
    new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_,
    new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_,
    new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_,
    new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_,
    new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_,
    new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_,
    new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_,
    new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_,
    new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6809_, new_n6810_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_,
    new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_,
    new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_,
    new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_,
    new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_,
    new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_,
    new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_,
    new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_,
    new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_,
    new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_,
    new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_,
    new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_,
    new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_,
    new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_,
    new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_,
    new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_,
    new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_,
    new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_,
    new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_,
    new_n6938_, new_n6939_, new_n6941_, new_n6942_, new_n6943_, new_n6944_,
    new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_,
    new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_,
    new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_,
    new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_,
    new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_,
    new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_,
    new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_,
    new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_,
    new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_,
    new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_,
    new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_,
    new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_,
    new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_,
    new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_,
    new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_,
    new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_,
    new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_,
    new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_,
    new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7058_, new_n7059_,
    new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_,
    new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_,
    new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_,
    new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_,
    new_n7084_, new_n7085_, new_n7086_, new_n7087_, new_n7088_, new_n7089_,
    new_n7090_, new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_,
    new_n7096_, new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_,
    new_n7102_, new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_,
    new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_,
    new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_,
    new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_,
    new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_, new_n7131_,
    new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_, new_n7137_,
    new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_, new_n7143_,
    new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_, new_n7149_,
    new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_, new_n7155_,
    new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_, new_n7161_,
    new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_, new_n7167_,
    new_n7168_, new_n7169_, new_n7170_, new_n7172_, new_n7173_, new_n7174_,
    new_n7175_, new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_,
    new_n7181_, new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_,
    new_n7187_, new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_,
    new_n7193_, new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_,
    new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_,
    new_n7205_, new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_,
    new_n7211_, new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_,
    new_n7217_, new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_,
    new_n7223_, new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_,
    new_n7229_, new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_,
    new_n7235_, new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_,
    new_n7241_, new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_,
    new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_,
    new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_,
    new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_, new_n7264_,
    new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_, new_n7270_,
    new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_, new_n7276_,
    new_n7277_, new_n7278_, new_n7279_, new_n7280_, new_n7281_, new_n7282_,
    new_n7283_, new_n7284_, new_n7286_, new_n7287_, new_n7288_, new_n7289_,
    new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_,
    new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_,
    new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_,
    new_n7308_, new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_,
    new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_,
    new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_,
    new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_,
    new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_,
    new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_,
    new_n7344_, new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_,
    new_n7350_, new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_,
    new_n7356_, new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_,
    new_n7362_, new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_,
    new_n7368_, new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_,
    new_n7374_, new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_,
    new_n7380_, new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_,
    new_n7386_, new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_,
    new_n7392_, new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_,
    new_n7398_, new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_,
    new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_,
    new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_,
    new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_,
    new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_,
    new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_,
    new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_,
    new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_,
    new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_,
    new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_,
    new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_,
    new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_,
    new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_,
    new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_,
    new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_,
    new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_,
    new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_,
    new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_,
    new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_,
    new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_,
    new_n7519_, new_n7520_, new_n7521_, new_n7523_, new_n7524_, new_n7525_,
    new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_,
    new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_,
    new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_,
    new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_,
    new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_,
    new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_,
    new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_,
    new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_,
    new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_,
    new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_,
    new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_,
    new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7639_, new_n7640_,
    new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_,
    new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_,
    new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_,
    new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_,
    new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_,
    new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_,
    new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_,
    new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_,
    new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_,
    new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_,
    new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_,
    new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_,
    new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_,
    new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_,
    new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_,
    new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_,
    new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_,
    new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_,
    new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_,
    new_n7755_, new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_,
    new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_,
    new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_,
    new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_,
    new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_,
    new_n7870_, new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_,
    new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_,
    new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_,
    new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_,
    new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_,
    new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_,
    new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_,
    new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_,
    new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_,
    new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_,
    new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_,
    new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7985_,
    new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_,
    new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_,
    new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_,
    new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_,
    new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8099_, new_n8100_,
    new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_,
    new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_,
    new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_,
    new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_,
    new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_,
    new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_,
    new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_,
    new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_,
    new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_,
    new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_,
    new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_,
    new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_,
    new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_,
    new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_,
    new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_,
    new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_,
    new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_,
    new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_,
    new_n8209_, new_n8210_, new_n8211_, new_n8213_, new_n8214_, new_n8215_,
    new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_,
    new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_,
    new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_,
    new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_,
    new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_, new_n8245_,
    new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_, new_n8251_,
    new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_,
    new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_, new_n8263_,
    new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_,
    new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_,
    new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_, new_n8281_,
    new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_,
    new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_, new_n8293_,
    new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_,
    new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_,
    new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_,
    new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_,
    new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_,
    new_n8324_, new_n8325_, new_n8326_, new_n8328_, new_n8329_, new_n8330_,
    new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_, new_n8336_,
    new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_, new_n8342_,
    new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_, new_n8348_,
    new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_, new_n8354_,
    new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_, new_n8360_,
    new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_, new_n8366_,
    new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8371_, new_n8372_,
    new_n8373_, new_n8374_, new_n8375_, new_n8376_, new_n8377_, new_n8378_,
    new_n8379_, new_n8380_, new_n8381_, new_n8382_, new_n8383_, new_n8384_,
    new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_, new_n8390_,
    new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_, new_n8396_,
    new_n8397_, new_n8398_, new_n8399_, new_n8400_, new_n8401_, new_n8402_,
    new_n8403_, new_n8404_, new_n8405_, new_n8406_, new_n8407_, new_n8408_,
    new_n8409_, new_n8410_, new_n8411_, new_n8412_, new_n8413_, new_n8414_,
    new_n8415_, new_n8416_, new_n8417_, new_n8418_, new_n8419_, new_n8420_,
    new_n8421_, new_n8422_, new_n8423_, new_n8424_, new_n8425_, new_n8426_,
    new_n8427_, new_n8428_, new_n8429_, new_n8430_, new_n8431_, new_n8432_,
    new_n8433_, new_n8434_, new_n8435_, new_n8436_, new_n8437_, new_n8438_,
    new_n8439_, new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_,
    new_n8446_, new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_,
    new_n8452_, new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_,
    new_n8458_, new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_,
    new_n8464_, new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_,
    new_n8470_, new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_,
    new_n8476_, new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_,
    new_n8482_, new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_,
    new_n8488_, new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_,
    new_n8494_, new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_,
    new_n8500_, new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_,
    new_n8506_, new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_,
    new_n8512_, new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_,
    new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_,
    new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8528_, new_n8529_,
    new_n8530_, new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_,
    new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_,
    new_n8542_, new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_,
    new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_,
    new_n8554_, new_n8555_, new_n8556_, new_n8557_, new_n8559_, new_n8560_,
    new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_,
    new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_,
    new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_,
    new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_,
    new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_,
    new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_,
    new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_,
    new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_,
    new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_,
    new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_,
    new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_,
    new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_,
    new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_,
    new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_,
    new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_,
    new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_,
    new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_,
    new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_,
    new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_,
    new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_,
    new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_,
    new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_,
    new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_,
    new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_,
    new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_,
    new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_,
    new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8789_, new_n8790_,
    new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_,
    new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_,
    new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_,
    new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_,
    new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_,
    new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_,
    new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_,
    new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_,
    new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_,
    new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_,
    new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_,
    new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_,
    new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_,
    new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_,
    new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_,
    new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_,
    new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_,
    new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_,
    new_n8899_, new_n8900_, new_n8901_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9023_, new_n9024_, new_n9025_, new_n9026_,
    new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_,
    new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_,
    new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_,
    new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_,
    new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_,
    new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_,
    new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_,
    new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_,
    new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_,
    new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_,
    new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_,
    new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_,
    new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_,
    new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_,
    new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_,
    new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_,
    new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_,
    new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_,
    new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9141_,
    new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_,
    new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_,
    new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_,
    new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_,
    new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_,
    new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_,
    new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_,
    new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_,
    new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_,
    new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_,
    new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_,
    new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_,
    new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_,
    new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_,
    new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_,
    new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_,
    new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_,
    new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_,
    new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_,
    new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_,
    new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_,
    new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_, new_n9274_,
    new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_, new_n9280_,
    new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_,
    new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_, new_n9292_,
    new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9298_,
    new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_, new_n9304_,
    new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_,
    new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_,
    new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_,
    new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_,
    new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_,
    new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_,
    new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_,
    new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_,
    new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_,
    new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_,
    new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_,
    new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_,
    new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_,
    new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_,
    new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_,
    new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_,
    new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_,
    new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_,
    new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_,
    new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_,
    new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_,
    new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_,
    new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_,
    new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_,
    new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_,
    new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_,
    new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_,
    new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_,
    new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_,
    new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_,
    new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_,
    new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_,
    new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_,
    new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_,
    new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_,
    new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_,
    new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_,
    new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_,
    new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_,
    new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_,
    new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_,
    new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_,
    new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_,
    new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_,
    new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_,
    new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_,
    new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_,
    new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_,
    new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_,
    new_n9601_, new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_,
    new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_,
    new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_,
    new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_,
    new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_,
    new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_, new_n9637_,
    new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_,
    new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_,
    new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_,
    new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_,
    new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_,
    new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_,
    new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_,
    new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_,
    new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_,
    new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_,
    new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_,
    new_n9716_, new_n9717_, new_n9719_, new_n9720_, new_n9721_, new_n9722_,
    new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_,
    new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_,
    new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_,
    new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_,
    new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_,
    new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_,
    new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_,
    new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_,
    new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_,
    new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_,
    new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_,
    new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_,
    new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_,
    new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_,
    new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_,
    new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_,
    new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_,
    new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9831_,
    new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_,
    new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_,
    new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_,
    new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_,
    new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_,
    new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_,
    new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_,
    new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_,
    new_n9881_, new_n9883_, new_n9885_, new_n9886_, new_n9887_, new_n9888_,
    new_n9889_, new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_,
    new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_,
    new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_,
    new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_,
    new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_,
    new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_,
    new_n9925_, new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_,
    new_n9931_, new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_,
    new_n9937_, new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_,
    new_n9943_, new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_,
    new_n9949_, new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_,
    new_n9955_, new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_,
    new_n9961_, new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_,
    new_n9967_, new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_,
    new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_,
    new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_,
    new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_,
    new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_,
    new_n9997_, new_n9998_, new_n10000_, new_n10001_, new_n10002_,
    new_n10003_, new_n10004_, new_n10005_, new_n10006_, new_n10007_,
    new_n10008_, new_n10009_, new_n10010_, new_n10011_, new_n10012_,
    new_n10013_, new_n10014_, new_n10015_, new_n10016_, new_n10017_,
    new_n10018_, new_n10019_, new_n10020_, new_n10021_, new_n10022_,
    new_n10023_, new_n10024_, new_n10025_, new_n10026_, new_n10027_,
    new_n10028_, new_n10029_, new_n10030_, new_n10031_, new_n10032_,
    new_n10033_, new_n10034_, new_n10035_, new_n10036_, new_n10037_,
    new_n10038_, new_n10039_, new_n10040_, new_n10041_, new_n10042_,
    new_n10043_, new_n10044_, new_n10045_, new_n10046_, new_n10047_,
    new_n10048_, new_n10049_, new_n10050_, new_n10051_, new_n10052_,
    new_n10053_, new_n10054_, new_n10055_, new_n10056_, new_n10057_,
    new_n10058_, new_n10059_, new_n10060_, new_n10061_, new_n10062_,
    new_n10063_, new_n10064_, new_n10065_, new_n10066_, new_n10067_,
    new_n10068_, new_n10069_, new_n10070_, new_n10071_, new_n10072_,
    new_n10073_, new_n10074_, new_n10075_, new_n10076_, new_n10077_,
    new_n10078_, new_n10079_, new_n10080_, new_n10081_, new_n10082_,
    new_n10083_, new_n10084_, new_n10085_, new_n10086_, new_n10087_,
    new_n10088_, new_n10089_, new_n10090_, new_n10091_, new_n10092_,
    new_n10093_, new_n10094_, new_n10095_, new_n10096_, new_n10097_,
    new_n10098_, new_n10099_, new_n10100_, new_n10101_, new_n10102_,
    new_n10103_, new_n10104_, new_n10105_, new_n10106_, new_n10107_,
    new_n10108_, new_n10109_, new_n10110_, new_n10111_, new_n10112_,
    new_n10113_, new_n10115_, new_n10116_, new_n10117_, new_n10118_,
    new_n10119_, new_n10120_, new_n10121_, new_n10122_, new_n10123_,
    new_n10124_, new_n10125_, new_n10126_, new_n10127_, new_n10128_,
    new_n10129_, new_n10130_, new_n10131_, new_n10132_, new_n10133_,
    new_n10134_, new_n10135_, new_n10136_, new_n10137_, new_n10138_,
    new_n10139_, new_n10140_, new_n10141_, new_n10142_, new_n10143_,
    new_n10144_, new_n10145_, new_n10146_, new_n10147_, new_n10148_,
    new_n10149_, new_n10150_, new_n10151_, new_n10152_, new_n10153_,
    new_n10154_, new_n10155_, new_n10156_, new_n10157_, new_n10158_,
    new_n10159_, new_n10160_, new_n10161_, new_n10162_, new_n10163_,
    new_n10164_, new_n10165_, new_n10166_, new_n10167_, new_n10168_,
    new_n10169_, new_n10170_, new_n10171_, new_n10172_, new_n10173_,
    new_n10174_, new_n10175_, new_n10176_, new_n10177_, new_n10178_,
    new_n10179_, new_n10180_, new_n10181_, new_n10182_, new_n10183_,
    new_n10184_, new_n10185_, new_n10186_, new_n10187_, new_n10188_,
    new_n10189_, new_n10190_, new_n10191_, new_n10192_, new_n10193_,
    new_n10194_, new_n10195_, new_n10196_, new_n10197_, new_n10198_,
    new_n10199_, new_n10200_, new_n10201_, new_n10202_, new_n10203_,
    new_n10204_, new_n10205_, new_n10206_, new_n10207_, new_n10208_,
    new_n10209_, new_n10210_, new_n10211_, new_n10212_, new_n10213_,
    new_n10214_, new_n10215_, new_n10216_, new_n10217_, new_n10218_,
    new_n10219_, new_n10220_, new_n10221_, new_n10222_, new_n10223_,
    new_n10224_, new_n10225_, new_n10226_, new_n10227_, new_n10228_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10460_, new_n10461_,
    new_n10462_, new_n10463_, new_n10464_, new_n10465_, new_n10466_,
    new_n10467_, new_n10468_, new_n10469_, new_n10470_, new_n10471_,
    new_n10472_, new_n10473_, new_n10474_, new_n10475_, new_n10476_,
    new_n10477_, new_n10478_, new_n10479_, new_n10480_, new_n10481_,
    new_n10482_, new_n10483_, new_n10484_, new_n10485_, new_n10486_,
    new_n10487_, new_n10488_, new_n10489_, new_n10490_, new_n10491_,
    new_n10492_, new_n10493_, new_n10494_, new_n10495_, new_n10496_,
    new_n10497_, new_n10498_, new_n10499_, new_n10500_, new_n10501_,
    new_n10502_, new_n10503_, new_n10504_, new_n10505_, new_n10506_,
    new_n10507_, new_n10508_, new_n10509_, new_n10510_, new_n10511_,
    new_n10512_, new_n10513_, new_n10514_, new_n10515_, new_n10516_,
    new_n10517_, new_n10518_, new_n10519_, new_n10520_, new_n10521_,
    new_n10522_, new_n10523_, new_n10524_, new_n10525_, new_n10526_,
    new_n10527_, new_n10528_, new_n10529_, new_n10530_, new_n10531_,
    new_n10532_, new_n10533_, new_n10534_, new_n10535_, new_n10536_,
    new_n10537_, new_n10538_, new_n10539_, new_n10540_, new_n10541_,
    new_n10542_, new_n10543_, new_n10544_, new_n10545_, new_n10546_,
    new_n10547_, new_n10548_, new_n10549_, new_n10550_, new_n10551_,
    new_n10552_, new_n10553_, new_n10554_, new_n10555_, new_n10556_,
    new_n10557_, new_n10558_, new_n10559_, new_n10560_, new_n10561_,
    new_n10562_, new_n10563_, new_n10564_, new_n10565_, new_n10566_,
    new_n10567_, new_n10568_, new_n10569_, new_n10570_, new_n10571_,
    new_n10572_, new_n10573_, new_n10574_, new_n10576_, new_n10577_,
    new_n10578_, new_n10579_, new_n10580_, new_n10581_, new_n10582_,
    new_n10583_, new_n10584_, new_n10585_, new_n10586_, new_n10587_,
    new_n10588_, new_n10589_, new_n10590_, new_n10591_, new_n10592_,
    new_n10593_, new_n10594_, new_n10595_, new_n10596_, new_n10597_,
    new_n10598_, new_n10599_, new_n10600_, new_n10601_, new_n10602_,
    new_n10603_, new_n10604_, new_n10605_, new_n10606_, new_n10607_,
    new_n10608_, new_n10609_, new_n10610_, new_n10611_, new_n10612_,
    new_n10613_, new_n10614_, new_n10615_, new_n10616_, new_n10617_,
    new_n10618_, new_n10619_, new_n10620_, new_n10621_, new_n10622_,
    new_n10623_, new_n10624_, new_n10625_, new_n10626_, new_n10627_,
    new_n10628_, new_n10629_, new_n10630_, new_n10631_, new_n10632_,
    new_n10633_, new_n10634_, new_n10635_, new_n10636_, new_n10637_,
    new_n10638_, new_n10639_, new_n10640_, new_n10641_, new_n10642_,
    new_n10643_, new_n10644_, new_n10645_, new_n10646_, new_n10647_,
    new_n10648_, new_n10649_, new_n10650_, new_n10651_, new_n10652_,
    new_n10653_, new_n10654_, new_n10655_, new_n10656_, new_n10657_,
    new_n10658_, new_n10659_, new_n10660_, new_n10661_, new_n10662_,
    new_n10663_, new_n10664_, new_n10665_, new_n10666_, new_n10667_,
    new_n10668_, new_n10669_, new_n10670_, new_n10671_, new_n10672_,
    new_n10673_, new_n10674_, new_n10675_, new_n10676_, new_n10677_,
    new_n10678_, new_n10679_, new_n10680_, new_n10681_, new_n10682_,
    new_n10683_, new_n10684_, new_n10685_, new_n10686_, new_n10687_,
    new_n10689_, new_n10690_, new_n10691_, new_n10692_, new_n10693_,
    new_n10694_, new_n10695_, new_n10696_, new_n10697_, new_n10698_,
    new_n10699_, new_n10700_, new_n10701_, new_n10702_, new_n10703_,
    new_n10704_, new_n10705_, new_n10706_, new_n10707_, new_n10708_,
    new_n10709_, new_n10710_, new_n10711_, new_n10712_, new_n10713_,
    new_n10714_, new_n10715_, new_n10716_, new_n10717_, new_n10718_,
    new_n10719_, new_n10720_, new_n10721_, new_n10722_, new_n10723_,
    new_n10724_, new_n10725_, new_n10726_, new_n10727_, new_n10728_,
    new_n10729_, new_n10730_, new_n10731_, new_n10732_, new_n10733_,
    new_n10734_, new_n10735_, new_n10736_, new_n10737_, new_n10738_,
    new_n10739_, new_n10740_, new_n10741_, new_n10742_, new_n10743_,
    new_n10744_, new_n10745_, new_n10746_, new_n10747_, new_n10748_,
    new_n10749_, new_n10750_, new_n10751_, new_n10752_, new_n10753_,
    new_n10754_, new_n10755_, new_n10756_, new_n10757_, new_n10758_,
    new_n10759_, new_n10760_, new_n10761_, new_n10762_, new_n10763_,
    new_n10764_, new_n10765_, new_n10766_, new_n10767_, new_n10768_,
    new_n10769_, new_n10770_, new_n10771_, new_n10772_, new_n10773_,
    new_n10774_, new_n10775_, new_n10776_, new_n10777_, new_n10778_,
    new_n10779_, new_n10780_, new_n10781_, new_n10782_, new_n10783_,
    new_n10784_, new_n10785_, new_n10786_, new_n10787_, new_n10788_,
    new_n10789_, new_n10790_, new_n10791_, new_n10792_, new_n10793_,
    new_n10794_, new_n10795_, new_n10796_, new_n10797_, new_n10798_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10817_, new_n10818_, new_n10819_,
    new_n10820_, new_n10821_, new_n10822_, new_n10823_, new_n10824_,
    new_n10825_, new_n10826_, new_n10827_, new_n10828_, new_n10829_,
    new_n10830_, new_n10831_, new_n10832_, new_n10833_, new_n10834_,
    new_n10835_, new_n10836_, new_n10837_, new_n10838_, new_n10839_,
    new_n10840_, new_n10841_, new_n10842_, new_n10843_, new_n10844_,
    new_n10845_, new_n10846_, new_n10847_, new_n10848_, new_n10849_,
    new_n10850_, new_n10851_, new_n10852_, new_n10853_, new_n10854_,
    new_n10855_, new_n10856_, new_n10857_, new_n10858_, new_n10859_,
    new_n10860_, new_n10861_, new_n10862_, new_n10863_, new_n10864_,
    new_n10865_, new_n10866_, new_n10867_, new_n10868_, new_n10869_,
    new_n10870_, new_n10871_, new_n10872_, new_n10873_, new_n10874_,
    new_n10875_, new_n10876_, new_n10877_, new_n10878_, new_n10879_,
    new_n10880_, new_n10881_, new_n10882_, new_n10883_, new_n10884_,
    new_n10885_, new_n10886_, new_n10887_, new_n10888_, new_n10889_,
    new_n10890_, new_n10891_, new_n10892_, new_n10893_, new_n10894_,
    new_n10895_, new_n10896_, new_n10897_, new_n10898_, new_n10899_,
    new_n10900_, new_n10901_, new_n10902_, new_n10903_, new_n10904_,
    new_n10905_, new_n10906_, new_n10907_, new_n10908_, new_n10909_,
    new_n10910_, new_n10911_, new_n10912_, new_n10913_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11030_, new_n11031_,
    new_n11032_, new_n11033_, new_n11034_, new_n11035_, new_n11036_,
    new_n11037_, new_n11038_, new_n11039_, new_n11040_, new_n11041_,
    new_n11042_, new_n11043_, new_n11044_, new_n11045_, new_n11046_,
    new_n11047_, new_n11048_, new_n11049_, new_n11050_, new_n11051_,
    new_n11052_, new_n11053_, new_n11054_, new_n11055_, new_n11056_,
    new_n11057_, new_n11058_, new_n11059_, new_n11060_, new_n11061_,
    new_n11062_, new_n11063_, new_n11064_, new_n11065_, new_n11066_,
    new_n11067_, new_n11068_, new_n11069_, new_n11070_, new_n11071_,
    new_n11072_, new_n11073_, new_n11074_, new_n11075_, new_n11076_,
    new_n11077_, new_n11078_, new_n11079_, new_n11080_, new_n11081_,
    new_n11082_, new_n11083_, new_n11084_, new_n11085_, new_n11086_,
    new_n11087_, new_n11088_, new_n11089_, new_n11090_, new_n11091_,
    new_n11092_, new_n11093_, new_n11094_, new_n11095_, new_n11096_,
    new_n11097_, new_n11098_, new_n11099_, new_n11100_, new_n11101_,
    new_n11102_, new_n11103_, new_n11104_, new_n11105_, new_n11106_,
    new_n11107_, new_n11108_, new_n11109_, new_n11110_, new_n11111_,
    new_n11112_, new_n11113_, new_n11114_, new_n11115_, new_n11116_,
    new_n11117_, new_n11118_, new_n11119_, new_n11120_, new_n11121_,
    new_n11122_, new_n11123_, new_n11124_, new_n11125_, new_n11126_,
    new_n11127_, new_n11128_, new_n11129_, new_n11130_, new_n11131_,
    new_n11132_, new_n11133_, new_n11134_, new_n11135_, new_n11136_,
    new_n11137_, new_n11138_, new_n11139_, new_n11140_, new_n11141_,
    new_n11142_, new_n11143_, new_n11144_, new_n11145_, new_n11147_,
    new_n11148_, new_n11149_, new_n11150_, new_n11151_, new_n11152_,
    new_n11153_, new_n11154_, new_n11155_, new_n11156_, new_n11157_,
    new_n11158_, new_n11159_, new_n11160_, new_n11161_, new_n11162_,
    new_n11163_, new_n11164_, new_n11165_, new_n11166_, new_n11167_,
    new_n11168_, new_n11169_, new_n11170_, new_n11171_, new_n11172_,
    new_n11173_, new_n11174_, new_n11175_, new_n11176_, new_n11177_,
    new_n11178_, new_n11179_, new_n11180_, new_n11181_, new_n11182_,
    new_n11183_, new_n11184_, new_n11185_, new_n11186_, new_n11187_,
    new_n11188_, new_n11189_, new_n11190_, new_n11191_, new_n11192_,
    new_n11193_, new_n11194_, new_n11195_, new_n11196_, new_n11197_,
    new_n11198_, new_n11199_, new_n11200_, new_n11201_, new_n11202_,
    new_n11203_, new_n11204_, new_n11205_, new_n11206_, new_n11207_,
    new_n11208_, new_n11209_, new_n11210_, new_n11211_, new_n11212_,
    new_n11213_, new_n11214_, new_n11215_, new_n11216_, new_n11217_,
    new_n11218_, new_n11219_, new_n11220_, new_n11221_, new_n11222_,
    new_n11223_, new_n11224_, new_n11225_, new_n11226_, new_n11227_,
    new_n11228_, new_n11229_, new_n11230_, new_n11231_, new_n11232_,
    new_n11233_, new_n11234_, new_n11235_, new_n11236_, new_n11237_,
    new_n11238_, new_n11239_, new_n11240_, new_n11241_, new_n11242_,
    new_n11243_, new_n11244_, new_n11245_, new_n11246_, new_n11247_,
    new_n11248_, new_n11249_, new_n11250_, new_n11251_, new_n11252_,
    new_n11253_, new_n11254_, new_n11255_, new_n11256_, new_n11257_,
    new_n11258_, new_n11259_, new_n11260_, new_n11261_, new_n11263_,
    new_n11264_, new_n11265_, new_n11266_, new_n11267_, new_n11268_,
    new_n11269_, new_n11270_, new_n11271_, new_n11272_, new_n11273_,
    new_n11274_, new_n11275_, new_n11276_, new_n11277_, new_n11278_,
    new_n11279_, new_n11280_, new_n11281_, new_n11282_, new_n11283_,
    new_n11284_, new_n11285_, new_n11286_, new_n11287_, new_n11288_,
    new_n11289_, new_n11290_, new_n11291_, new_n11292_, new_n11293_,
    new_n11294_, new_n11295_, new_n11296_, new_n11297_, new_n11298_,
    new_n11299_, new_n11300_, new_n11301_, new_n11302_, new_n11303_,
    new_n11304_, new_n11305_, new_n11306_, new_n11307_, new_n11308_,
    new_n11309_, new_n11310_, new_n11311_, new_n11312_, new_n11313_,
    new_n11314_, new_n11315_, new_n11316_, new_n11317_, new_n11318_,
    new_n11319_, new_n11320_, new_n11321_, new_n11322_, new_n11323_,
    new_n11324_, new_n11325_, new_n11326_, new_n11327_, new_n11328_,
    new_n11329_, new_n11330_, new_n11331_, new_n11332_, new_n11333_,
    new_n11334_, new_n11335_, new_n11336_, new_n11337_, new_n11338_,
    new_n11339_, new_n11340_, new_n11341_, new_n11342_, new_n11343_,
    new_n11344_, new_n11345_, new_n11346_, new_n11347_, new_n11348_,
    new_n11349_, new_n11350_, new_n11351_, new_n11352_, new_n11353_,
    new_n11354_, new_n11355_, new_n11356_, new_n11357_, new_n11358_,
    new_n11359_, new_n11360_, new_n11361_, new_n11362_, new_n11363_,
    new_n11364_, new_n11365_, new_n11366_, new_n11367_, new_n11368_,
    new_n11369_, new_n11370_, new_n11371_, new_n11372_, new_n11373_,
    new_n11374_, new_n11375_, new_n11376_, new_n11378_, new_n11379_,
    new_n11380_, new_n11381_, new_n11382_, new_n11383_, new_n11384_,
    new_n11385_, new_n11386_, new_n11387_, new_n11388_, new_n11389_,
    new_n11390_, new_n11391_, new_n11392_, new_n11393_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11399_,
    new_n11400_, new_n11401_, new_n11402_, new_n11403_, new_n11404_,
    new_n11405_, new_n11406_, new_n11407_, new_n11408_, new_n11409_,
    new_n11410_, new_n11411_, new_n11412_, new_n11413_, new_n11414_,
    new_n11415_, new_n11416_, new_n11417_, new_n11418_, new_n11419_,
    new_n11420_, new_n11421_, new_n11422_, new_n11423_, new_n11424_,
    new_n11425_, new_n11426_, new_n11427_, new_n11428_, new_n11429_,
    new_n11430_, new_n11431_, new_n11432_, new_n11433_, new_n11434_,
    new_n11435_, new_n11436_, new_n11437_, new_n11438_, new_n11439_,
    new_n11440_, new_n11441_, new_n11442_, new_n11443_, new_n11444_,
    new_n11445_, new_n11446_, new_n11447_, new_n11448_, new_n11449_,
    new_n11450_, new_n11451_, new_n11452_, new_n11453_, new_n11454_,
    new_n11455_, new_n11456_, new_n11457_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11491_, new_n11492_, new_n11493_, new_n11494_, new_n11495_,
    new_n11496_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11503_, new_n11504_, new_n11505_,
    new_n11506_, new_n11507_, new_n11508_, new_n11509_, new_n11510_,
    new_n11511_, new_n11512_, new_n11513_, new_n11514_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11618_, new_n11619_, new_n11620_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11645_, new_n11646_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11652_, new_n11653_, new_n11654_, new_n11655_, new_n11656_,
    new_n11657_, new_n11658_, new_n11659_, new_n11660_, new_n11661_,
    new_n11662_, new_n11663_, new_n11664_, new_n11665_, new_n11666_,
    new_n11667_, new_n11668_, new_n11669_, new_n11670_, new_n11671_,
    new_n11672_, new_n11673_, new_n11674_, new_n11675_, new_n11676_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11682_, new_n11683_, new_n11684_, new_n11685_, new_n11686_,
    new_n11687_, new_n11688_, new_n11689_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11712_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11721_,
    new_n11722_, new_n11723_, new_n11724_, new_n11725_, new_n11726_,
    new_n11727_, new_n11729_, new_n11730_, new_n11731_, new_n11732_,
    new_n11733_, new_n11734_, new_n11735_, new_n11736_, new_n11737_,
    new_n11738_, new_n11739_, new_n11740_, new_n11741_, new_n11742_,
    new_n11743_, new_n11744_, new_n11745_, new_n11746_, new_n11747_,
    new_n11748_, new_n11749_, new_n11750_, new_n11751_, new_n11752_,
    new_n11753_, new_n11754_, new_n11755_, new_n11756_, new_n11757_,
    new_n11758_, new_n11759_, new_n11760_, new_n11761_, new_n11762_,
    new_n11763_, new_n11764_, new_n11765_, new_n11766_, new_n11767_,
    new_n11768_, new_n11769_, new_n11770_, new_n11771_, new_n11772_,
    new_n11773_, new_n11774_, new_n11775_, new_n11776_, new_n11777_,
    new_n11778_, new_n11779_, new_n11780_, new_n11781_, new_n11782_,
    new_n11783_, new_n11784_, new_n11785_, new_n11786_, new_n11787_,
    new_n11788_, new_n11789_, new_n11790_, new_n11791_, new_n11792_,
    new_n11793_, new_n11794_, new_n11795_, new_n11796_, new_n11797_,
    new_n11798_, new_n11799_, new_n11800_, new_n11801_, new_n11802_,
    new_n11803_, new_n11804_, new_n11805_, new_n11806_, new_n11807_,
    new_n11808_, new_n11809_, new_n11810_, new_n11811_, new_n11812_,
    new_n11813_, new_n11814_, new_n11815_, new_n11816_, new_n11817_,
    new_n11818_, new_n11819_, new_n11820_, new_n11821_, new_n11822_,
    new_n11823_, new_n11824_, new_n11825_, new_n11826_, new_n11827_,
    new_n11828_, new_n11829_, new_n11830_, new_n11831_, new_n11832_,
    new_n11833_, new_n11834_, new_n11835_, new_n11836_, new_n11837_,
    new_n11838_, new_n11839_, new_n11840_, new_n11841_, new_n11842_,
    new_n11843_, new_n11845_, new_n11846_, new_n11847_, new_n11848_,
    new_n11849_, new_n11850_, new_n11851_, new_n11852_, new_n11853_,
    new_n11854_, new_n11855_, new_n11856_, new_n11857_, new_n11858_,
    new_n11859_, new_n11860_, new_n11861_, new_n11862_, new_n11863_,
    new_n11864_, new_n11865_, new_n11866_, new_n11867_, new_n11868_,
    new_n11869_, new_n11870_, new_n11871_, new_n11872_, new_n11873_,
    new_n11874_, new_n11875_, new_n11876_, new_n11877_, new_n11878_,
    new_n11879_, new_n11880_, new_n11881_, new_n11882_, new_n11883_,
    new_n11884_, new_n11885_, new_n11886_, new_n11887_, new_n11888_,
    new_n11889_, new_n11890_, new_n11891_, new_n11892_, new_n11893_,
    new_n11894_, new_n11895_, new_n11896_, new_n11897_, new_n11898_,
    new_n11899_, new_n11900_, new_n11901_, new_n11902_, new_n11903_,
    new_n11904_, new_n11905_, new_n11906_, new_n11907_, new_n11908_,
    new_n11909_, new_n11910_, new_n11911_, new_n11912_, new_n11913_,
    new_n11914_, new_n11915_, new_n11916_, new_n11917_, new_n11918_,
    new_n11919_, new_n11920_, new_n11921_, new_n11922_, new_n11923_,
    new_n11924_, new_n11925_, new_n11926_, new_n11927_, new_n11928_,
    new_n11929_, new_n11930_, new_n11931_, new_n11932_, new_n11933_,
    new_n11934_, new_n11935_, new_n11936_, new_n11937_, new_n11938_,
    new_n11939_, new_n11940_, new_n11941_, new_n11942_, new_n11943_,
    new_n11944_, new_n11945_, new_n11946_, new_n11947_, new_n11948_,
    new_n11949_, new_n11950_, new_n11951_, new_n11952_, new_n11953_,
    new_n11954_, new_n11955_, new_n11956_, new_n11957_, new_n11958_,
    new_n11959_, new_n11961_, new_n11962_, new_n11963_, new_n11964_,
    new_n11965_, new_n11966_, new_n11967_, new_n11968_, new_n11969_,
    new_n11970_, new_n11972_, new_n11973_, new_n11974_, new_n11975_,
    new_n11976_, new_n11977_, new_n11978_, new_n11979_, new_n11980_,
    new_n11981_, new_n11982_, new_n11983_, new_n11984_, new_n11985_,
    new_n11986_, new_n11987_, new_n11988_, new_n11989_, new_n11990_,
    new_n11991_, new_n11992_, new_n11993_, new_n11994_, new_n11995_,
    new_n11996_, new_n11997_, new_n11998_, new_n11999_, new_n12000_,
    new_n12001_, new_n12002_, new_n12003_, new_n12004_, new_n12005_,
    new_n12006_, new_n12007_, new_n12008_, new_n12009_, new_n12010_,
    new_n12011_, new_n12012_, new_n12013_, new_n12014_, new_n12015_,
    new_n12016_, new_n12017_, new_n12018_, new_n12019_, new_n12020_,
    new_n12021_, new_n12022_, new_n12023_, new_n12024_, new_n12025_,
    new_n12026_, new_n12027_, new_n12028_, new_n12029_, new_n12030_,
    new_n12031_, new_n12032_, new_n12033_, new_n12034_, new_n12035_,
    new_n12036_, new_n12037_, new_n12038_, new_n12039_, new_n12040_,
    new_n12041_, new_n12042_, new_n12043_, new_n12044_, new_n12045_,
    new_n12046_, new_n12047_, new_n12048_, new_n12049_, new_n12050_,
    new_n12051_, new_n12052_, new_n12053_, new_n12054_, new_n12055_,
    new_n12056_, new_n12057_, new_n12058_, new_n12059_, new_n12060_,
    new_n12061_, new_n12062_, new_n12063_, new_n12064_, new_n12065_,
    new_n12066_, new_n12067_, new_n12068_, new_n12069_, new_n12070_,
    new_n12071_, new_n12072_, new_n12073_, new_n12074_, new_n12075_,
    new_n12076_, new_n12077_, new_n12078_, new_n12079_, new_n12080_,
    new_n12081_, new_n12082_, new_n12083_, new_n12084_, new_n12085_,
    new_n12086_, new_n12088_, new_n12089_, new_n12090_, new_n12091_,
    new_n12092_, new_n12093_, new_n12094_, new_n12096_, new_n12097_,
    new_n12098_, new_n12099_, new_n12100_, new_n12101_, new_n12102_,
    new_n12103_, new_n12104_, new_n12105_, new_n12106_, new_n12107_,
    new_n12108_, new_n12109_, new_n12110_, new_n12111_, new_n12112_,
    new_n12113_, new_n12114_, new_n12115_, new_n12116_, new_n12117_,
    new_n12118_, new_n12119_, new_n12120_, new_n12121_, new_n12122_,
    new_n12123_, new_n12124_, new_n12125_, new_n12126_, new_n12127_,
    new_n12128_, new_n12129_, new_n12130_, new_n12131_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12136_, new_n12137_,
    new_n12138_, new_n12139_, new_n12140_, new_n12141_, new_n12142_,
    new_n12143_, new_n12144_, new_n12145_, new_n12146_, new_n12147_,
    new_n12148_, new_n12149_, new_n12150_, new_n12151_, new_n12152_,
    new_n12153_, new_n12154_, new_n12155_, new_n12156_, new_n12157_,
    new_n12158_, new_n12159_, new_n12160_, new_n12161_, new_n12162_,
    new_n12163_, new_n12164_, new_n12165_, new_n12166_, new_n12167_,
    new_n12168_, new_n12169_, new_n12170_, new_n12171_, new_n12172_,
    new_n12173_, new_n12174_, new_n12175_, new_n12176_, new_n12177_,
    new_n12178_, new_n12179_, new_n12180_, new_n12181_, new_n12182_,
    new_n12183_, new_n12184_, new_n12185_, new_n12186_, new_n12187_,
    new_n12188_, new_n12189_, new_n12190_, new_n12191_, new_n12192_,
    new_n12193_, new_n12194_, new_n12195_, new_n12196_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12203_, new_n12204_, new_n12205_, new_n12206_, new_n12207_,
    new_n12208_, new_n12210_, new_n12211_, new_n12212_, new_n12213_,
    new_n12214_, new_n12215_, new_n12216_, new_n12217_, new_n12218_,
    new_n12219_, new_n12220_, new_n12221_, new_n12222_, new_n12223_,
    new_n12224_, new_n12225_, new_n12226_, new_n12227_, new_n12228_,
    new_n12229_, new_n12230_, new_n12231_, new_n12232_, new_n12233_,
    new_n12234_, new_n12235_, new_n12236_, new_n12237_, new_n12238_,
    new_n12239_, new_n12240_, new_n12241_, new_n12242_, new_n12243_,
    new_n12244_, new_n12245_, new_n12246_, new_n12247_, new_n12248_,
    new_n12249_, new_n12250_, new_n12251_, new_n12252_, new_n12253_,
    new_n12254_, new_n12255_, new_n12256_, new_n12257_, new_n12258_,
    new_n12259_, new_n12260_, new_n12261_, new_n12262_, new_n12263_,
    new_n12264_, new_n12265_, new_n12266_, new_n12267_, new_n12268_,
    new_n12269_, new_n12270_, new_n12271_, new_n12272_, new_n12273_,
    new_n12274_, new_n12275_, new_n12276_, new_n12277_, new_n12278_,
    new_n12279_, new_n12280_, new_n12281_, new_n12282_, new_n12283_,
    new_n12284_, new_n12285_, new_n12286_, new_n12287_, new_n12288_,
    new_n12289_, new_n12290_, new_n12291_, new_n12292_, new_n12293_,
    new_n12294_, new_n12295_, new_n12296_, new_n12297_, new_n12298_,
    new_n12299_, new_n12300_, new_n12301_, new_n12302_, new_n12303_,
    new_n12304_, new_n12305_, new_n12306_, new_n12307_, new_n12308_,
    new_n12309_, new_n12310_, new_n12311_, new_n12312_, new_n12313_,
    new_n12314_, new_n12315_, new_n12316_, new_n12317_, new_n12318_,
    new_n12319_, new_n12320_, new_n12321_, new_n12322_, new_n12324_,
    new_n12325_, new_n12326_, new_n12327_, new_n12328_, new_n12329_,
    new_n12330_, new_n12331_, new_n12332_, new_n12333_, new_n12334_,
    new_n12335_, new_n12336_, new_n12337_, new_n12338_, new_n12339_,
    new_n12340_, new_n12341_, new_n12342_, new_n12343_, new_n12344_,
    new_n12345_, new_n12346_, new_n12347_, new_n12348_, new_n12349_,
    new_n12350_, new_n12351_, new_n12352_, new_n12353_, new_n12354_,
    new_n12355_, new_n12356_, new_n12357_, new_n12358_, new_n12359_,
    new_n12360_, new_n12361_, new_n12362_, new_n12363_, new_n12364_,
    new_n12365_, new_n12366_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12375_, new_n12376_, new_n12377_, new_n12378_, new_n12379_,
    new_n12380_, new_n12381_, new_n12382_, new_n12383_, new_n12384_,
    new_n12385_, new_n12386_, new_n12387_, new_n12388_, new_n12389_,
    new_n12390_, new_n12391_, new_n12392_, new_n12393_, new_n12394_,
    new_n12395_, new_n12396_, new_n12397_, new_n12398_, new_n12399_,
    new_n12400_, new_n12401_, new_n12402_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12409_,
    new_n12410_, new_n12411_, new_n12412_, new_n12413_, new_n12414_,
    new_n12415_, new_n12416_, new_n12417_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12438_, new_n12439_, new_n12440_,
    new_n12441_, new_n12442_, new_n12443_, new_n12444_, new_n12445_,
    new_n12446_, new_n12447_, new_n12448_, new_n12449_, new_n12450_,
    new_n12451_, new_n12452_, new_n12453_, new_n12454_, new_n12455_,
    new_n12456_, new_n12457_, new_n12458_, new_n12459_, new_n12460_,
    new_n12461_, new_n12462_, new_n12463_, new_n12464_, new_n12465_,
    new_n12466_, new_n12467_, new_n12468_, new_n12469_, new_n12470_,
    new_n12471_, new_n12472_, new_n12473_, new_n12474_, new_n12475_,
    new_n12476_, new_n12477_, new_n12478_, new_n12479_, new_n12480_,
    new_n12481_, new_n12482_, new_n12483_, new_n12484_, new_n12485_,
    new_n12486_, new_n12487_, new_n12488_, new_n12489_, new_n12490_,
    new_n12491_, new_n12492_, new_n12493_, new_n12494_, new_n12495_,
    new_n12496_, new_n12497_, new_n12498_, new_n12499_, new_n12500_,
    new_n12501_, new_n12502_, new_n12503_, new_n12504_, new_n12505_,
    new_n12506_, new_n12507_, new_n12508_, new_n12509_, new_n12510_,
    new_n12511_, new_n12512_, new_n12513_, new_n12514_, new_n12515_,
    new_n12516_, new_n12517_, new_n12518_, new_n12519_, new_n12520_,
    new_n12521_, new_n12522_, new_n12523_, new_n12524_, new_n12525_,
    new_n12526_, new_n12527_, new_n12528_, new_n12529_, new_n12530_,
    new_n12531_, new_n12532_, new_n12533_, new_n12534_, new_n12535_,
    new_n12536_, new_n12537_, new_n12538_, new_n12539_, new_n12540_,
    new_n12541_, new_n12542_, new_n12543_, new_n12544_, new_n12545_,
    new_n12546_, new_n12547_, new_n12548_, new_n12549_, new_n12550_,
    new_n12552_, new_n12553_, new_n12554_, new_n12555_, new_n12556_,
    new_n12557_, new_n12558_, new_n12559_, new_n12560_, new_n12561_,
    new_n12562_, new_n12563_, new_n12564_, new_n12565_, new_n12566_,
    new_n12567_, new_n12568_, new_n12569_, new_n12570_, new_n12571_,
    new_n12572_, new_n12573_, new_n12574_, new_n12575_, new_n12576_,
    new_n12577_, new_n12578_, new_n12579_, new_n12580_, new_n12581_,
    new_n12582_, new_n12583_, new_n12584_, new_n12585_, new_n12586_,
    new_n12587_, new_n12588_, new_n12589_, new_n12590_, new_n12591_,
    new_n12592_, new_n12593_, new_n12594_, new_n12595_, new_n12596_,
    new_n12597_, new_n12598_, new_n12599_, new_n12600_, new_n12601_,
    new_n12602_, new_n12603_, new_n12604_, new_n12605_, new_n12606_,
    new_n12607_, new_n12608_, new_n12609_, new_n12610_, new_n12611_,
    new_n12612_, new_n12613_, new_n12614_, new_n12615_, new_n12616_,
    new_n12617_, new_n12618_, new_n12619_, new_n12620_, new_n12621_,
    new_n12622_, new_n12623_, new_n12624_, new_n12625_, new_n12626_,
    new_n12627_, new_n12628_, new_n12629_, new_n12630_, new_n12631_,
    new_n12632_, new_n12633_, new_n12634_, new_n12635_, new_n12636_,
    new_n12637_, new_n12638_, new_n12639_, new_n12640_, new_n12641_,
    new_n12642_, new_n12643_, new_n12644_, new_n12645_, new_n12646_,
    new_n12647_, new_n12648_, new_n12649_, new_n12650_, new_n12651_,
    new_n12652_, new_n12653_, new_n12654_, new_n12655_, new_n12656_,
    new_n12657_, new_n12658_, new_n12659_, new_n12660_, new_n12661_,
    new_n12662_, new_n12663_, new_n12665_, new_n12666_, new_n12667_,
    new_n12668_, new_n12669_, new_n12670_, new_n12671_, new_n12672_,
    new_n12673_, new_n12674_, new_n12675_, new_n12676_, new_n12677_,
    new_n12678_, new_n12679_, new_n12680_, new_n12681_, new_n12682_,
    new_n12683_, new_n12684_, new_n12685_, new_n12686_, new_n12687_,
    new_n12688_, new_n12689_, new_n12690_, new_n12691_, new_n12692_,
    new_n12693_, new_n12694_, new_n12695_, new_n12696_, new_n12697_,
    new_n12698_, new_n12699_, new_n12700_, new_n12701_, new_n12702_,
    new_n12703_, new_n12704_, new_n12705_, new_n12706_, new_n12707_,
    new_n12708_, new_n12709_, new_n12710_, new_n12711_, new_n12712_,
    new_n12713_, new_n12714_, new_n12715_, new_n12716_, new_n12717_,
    new_n12718_, new_n12719_, new_n12720_, new_n12721_, new_n12722_,
    new_n12723_, new_n12724_, new_n12725_, new_n12726_, new_n12727_,
    new_n12728_, new_n12729_, new_n12730_, new_n12731_, new_n12732_,
    new_n12733_, new_n12734_, new_n12735_, new_n12736_, new_n12737_,
    new_n12738_, new_n12739_, new_n12740_, new_n12741_, new_n12742_,
    new_n12743_, new_n12744_, new_n12745_, new_n12746_, new_n12747_,
    new_n12748_, new_n12749_, new_n12750_, new_n12751_, new_n12752_,
    new_n12753_, new_n12754_, new_n12755_, new_n12756_, new_n12757_,
    new_n12758_, new_n12759_, new_n12760_, new_n12761_, new_n12762_,
    new_n12763_, new_n12764_, new_n12765_, new_n12766_, new_n12767_,
    new_n12768_, new_n12769_, new_n12770_, new_n12771_, new_n12772_,
    new_n12773_, new_n12774_, new_n12775_, new_n12776_, new_n12777_,
    new_n12778_, new_n12779_, new_n12781_, new_n12782_, new_n12783_,
    new_n12784_, new_n12785_, new_n12786_, new_n12787_, new_n12788_,
    new_n12789_, new_n12790_, new_n12791_, new_n12792_, new_n12793_,
    new_n12794_, new_n12795_, new_n12796_, new_n12797_, new_n12798_,
    new_n12799_, new_n12800_, new_n12801_, new_n12802_, new_n12803_,
    new_n12804_, new_n12805_, new_n12806_, new_n12807_, new_n12808_,
    new_n12809_, new_n12810_, new_n12811_, new_n12812_, new_n12813_,
    new_n12814_, new_n12815_, new_n12816_, new_n12817_, new_n12818_,
    new_n12819_, new_n12820_, new_n12821_, new_n12822_, new_n12823_,
    new_n12824_, new_n12825_, new_n12826_, new_n12827_, new_n12828_,
    new_n12829_, new_n12830_, new_n12831_, new_n12832_, new_n12833_,
    new_n12834_, new_n12835_, new_n12836_, new_n12837_, new_n12838_,
    new_n12839_, new_n12840_, new_n12841_, new_n12842_, new_n12843_,
    new_n12844_, new_n12845_, new_n12846_, new_n12847_, new_n12848_,
    new_n12849_, new_n12850_, new_n12851_, new_n12852_, new_n12853_,
    new_n12854_, new_n12855_, new_n12856_, new_n12857_, new_n12858_,
    new_n12859_, new_n12860_, new_n12861_, new_n12862_, new_n12863_,
    new_n12864_, new_n12865_, new_n12866_, new_n12867_, new_n12868_,
    new_n12869_, new_n12870_, new_n12871_, new_n12872_, new_n12873_,
    new_n12874_, new_n12875_, new_n12876_, new_n12877_, new_n12878_,
    new_n12879_, new_n12880_, new_n12881_, new_n12882_, new_n12883_,
    new_n12884_, new_n12885_, new_n12886_, new_n12887_, new_n12888_,
    new_n12889_, new_n12890_, new_n12891_, new_n12892_, new_n12893_,
    new_n12894_, new_n12895_, new_n12897_, new_n12898_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13006_, new_n13007_, new_n13008_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13126_, new_n13127_,
    new_n13128_, new_n13129_, new_n13130_, new_n13131_, new_n13133_,
    new_n13134_, new_n13135_, new_n13136_, new_n13137_, new_n13138_,
    new_n13139_, new_n13141_, new_n13142_, new_n13143_, new_n13144_,
    new_n13145_, new_n13146_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13155_, new_n13156_,
    new_n13157_, new_n13158_, new_n13159_, new_n13160_, new_n13161_,
    new_n13163_, new_n13164_, new_n13165_, new_n13166_, new_n13167_,
    new_n13168_, new_n13169_, new_n13170_, new_n13171_, new_n13172_,
    new_n13173_, new_n13174_, new_n13175_, new_n13176_, new_n13177_,
    new_n13178_, new_n13179_, new_n13180_, new_n13181_, new_n13182_,
    new_n13183_, new_n13184_, new_n13185_, new_n13186_, new_n13187_,
    new_n13188_, new_n13189_, new_n13190_, new_n13191_, new_n13192_,
    new_n13193_, new_n13194_, new_n13195_, new_n13196_, new_n13197_,
    new_n13198_, new_n13199_, new_n13200_, new_n13201_, new_n13202_,
    new_n13203_, new_n13205_, new_n13206_, new_n13207_, new_n13208_,
    new_n13209_, new_n13210_, new_n13211_, new_n13212_, new_n13213_,
    new_n13214_, new_n13215_, new_n13216_, new_n13217_, new_n13219_,
    new_n13220_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13228_, new_n13229_, new_n13231_, new_n13232_,
    new_n13233_, new_n13234_, new_n13235_, new_n13236_, new_n13237_,
    new_n13238_, new_n13239_, new_n13240_, new_n13241_, new_n13242_,
    new_n13243_, new_n13244_, new_n13245_, new_n13246_, new_n13247_,
    new_n13248_, new_n13249_, new_n13250_, new_n13251_, new_n13252_,
    new_n13253_, new_n13254_, new_n13255_, new_n13256_, new_n13257_,
    new_n13258_, new_n13259_, new_n13260_, new_n13261_, new_n13262_,
    new_n13263_, new_n13264_, new_n13265_, new_n13266_, new_n13267_,
    new_n13268_, new_n13269_, new_n13270_, new_n13271_, new_n13272_,
    new_n13273_, new_n13274_, new_n13275_, new_n13277_, new_n13278_,
    new_n13279_, new_n13280_, new_n13281_, new_n13282_, new_n13283_,
    new_n13284_, new_n13285_, new_n13286_, new_n13287_, new_n13288_,
    new_n13289_, new_n13290_, new_n13291_, new_n13292_, new_n13293_,
    new_n13294_, new_n13295_, new_n13296_, new_n13297_, new_n13298_,
    new_n13299_, new_n13300_, new_n13301_, new_n13302_, new_n13303_,
    new_n13304_, new_n13305_, new_n13306_, new_n13307_, new_n13308_,
    new_n13309_, new_n13310_, new_n13311_, new_n13312_, new_n13313_,
    new_n13314_, new_n13315_, new_n13316_, new_n13317_, new_n13318_,
    new_n13319_, new_n13320_, new_n13321_, new_n13322_, new_n13323_,
    new_n13324_, new_n13325_, new_n13326_, new_n13327_, new_n13328_,
    new_n13329_, new_n13330_, new_n13331_, new_n13332_, new_n13333_,
    new_n13334_, new_n13335_, new_n13336_, new_n13337_, new_n13338_,
    new_n13339_, new_n13340_, new_n13341_, new_n13342_, new_n13343_,
    new_n13344_, new_n13345_, new_n13346_, new_n13347_, new_n13348_,
    new_n13349_, new_n13350_, new_n13351_, new_n13352_, new_n13353_,
    new_n13354_, new_n13355_, new_n13356_, new_n13357_, new_n13358_,
    new_n13359_, new_n13360_, new_n13361_, new_n13362_, new_n13363_,
    new_n13364_, new_n13365_, new_n13366_, new_n13367_, new_n13368_,
    new_n13369_, new_n13370_, new_n13371_, new_n13372_, new_n13373_,
    new_n13374_, new_n13375_, new_n13376_, new_n13377_, new_n13378_,
    new_n13379_, new_n13380_, new_n13381_, new_n13382_, new_n13384_,
    new_n13385_, new_n13386_, new_n13387_, new_n13388_, new_n13389_,
    new_n13390_, new_n13391_, new_n13392_, new_n13393_, new_n13394_,
    new_n13395_, new_n13396_, new_n13397_, new_n13398_, new_n13399_,
    new_n13400_, new_n13401_, new_n13402_, new_n13403_, new_n13404_,
    new_n13405_, new_n13406_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13435_, new_n13436_,
    new_n13437_, new_n13438_, new_n13439_, new_n13440_, new_n13441_,
    new_n13442_, new_n13443_, new_n13444_, new_n13445_, new_n13446_,
    new_n13447_, new_n13448_, new_n13449_, new_n13450_, new_n13451_,
    new_n13452_, new_n13453_, new_n13454_, new_n13455_, new_n13456_,
    new_n13457_, new_n13458_, new_n13459_, new_n13460_, new_n13461_,
    new_n13462_, new_n13463_, new_n13464_, new_n13465_, new_n13466_,
    new_n13467_, new_n13468_, new_n13469_, new_n13470_, new_n13471_,
    new_n13472_, new_n13474_, new_n13475_, new_n13476_, new_n13477_,
    new_n13478_, new_n13479_, new_n13480_, new_n13481_, new_n13482_,
    new_n13483_, new_n13484_, new_n13485_, new_n13486_, new_n13487_,
    new_n13488_, new_n13489_, new_n13490_, new_n13491_, new_n13492_,
    new_n13493_, new_n13494_, new_n13496_, new_n13497_, new_n13498_,
    new_n13499_, new_n13500_, new_n13501_, new_n13502_, new_n13503_,
    new_n13504_, new_n13505_, new_n13506_, new_n13507_, new_n13508_,
    new_n13509_, new_n13510_, new_n13511_, new_n13513_, new_n13514_,
    new_n13515_, new_n13516_, new_n13517_, new_n13518_, new_n13519_,
    new_n13520_, new_n13521_, new_n13522_, new_n13523_, new_n13524_,
    new_n13525_, new_n13526_, new_n13527_, new_n13528_, new_n13529_,
    new_n13530_, new_n13531_, new_n13532_, new_n13533_, new_n13534_,
    new_n13535_, new_n13536_, new_n13537_, new_n13538_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13575_, new_n13576_, new_n13577_,
    new_n13578_, new_n13579_, new_n13580_, new_n13581_, new_n13582_,
    new_n13583_, new_n13584_, new_n13585_, new_n13586_, new_n13587_,
    new_n13588_, new_n13589_, new_n13590_, new_n13591_, new_n13593_,
    new_n13594_, new_n13595_, new_n13596_, new_n13597_, new_n13598_,
    new_n13599_, new_n13600_, new_n13601_, new_n13602_, new_n13603_,
    new_n13604_, new_n13605_, new_n13606_, new_n13607_, new_n13608_,
    new_n13610_, new_n13611_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13620_,
    new_n13621_, new_n13622_, new_n13623_, new_n13624_, new_n13625_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13638_, new_n13639_, new_n13640_, new_n13641_, new_n13642_,
    new_n13643_, new_n13644_, new_n13645_, new_n13646_, new_n13647_,
    new_n13648_, new_n13649_, new_n13650_, new_n13651_, new_n13652_,
    new_n13653_, new_n13654_, new_n13655_, new_n13656_, new_n13657_,
    new_n13658_, new_n13659_, new_n13660_, new_n13661_, new_n13662_,
    new_n13663_, new_n13664_, new_n13665_, new_n13666_, new_n13668_,
    new_n13669_, new_n13670_, new_n13671_, new_n13672_, new_n13673_,
    new_n13674_, new_n13675_, new_n13676_, new_n13677_, new_n13678_,
    new_n13679_, new_n13680_, new_n13681_, new_n13682_, new_n13683_,
    new_n13684_, new_n13685_, new_n13686_, new_n13687_, new_n13688_,
    new_n13689_, new_n13690_, new_n13691_, new_n13692_, new_n13693_,
    new_n13694_, new_n13695_, new_n13696_, new_n13697_, new_n13698_,
    new_n13699_, new_n13700_, new_n13701_, new_n13702_, new_n13703_,
    new_n13704_, new_n13705_, new_n13706_, new_n13707_, new_n13708_,
    new_n13709_, new_n13710_, new_n13711_, new_n13712_, new_n13713_,
    new_n13714_, new_n13715_, new_n13716_, new_n13717_, new_n13718_,
    new_n13719_, new_n13720_, new_n13721_, new_n13722_, new_n13723_,
    new_n13724_, new_n13725_, new_n13726_, new_n13727_, new_n13728_,
    new_n13729_, new_n13730_, new_n13731_, new_n13732_, new_n13733_,
    new_n13734_, new_n13735_, new_n13736_, new_n13737_, new_n13738_,
    new_n13739_, new_n13740_, new_n13741_, new_n13742_, new_n13743_,
    new_n13744_, new_n13745_, new_n13746_, new_n13747_, new_n13748_,
    new_n13749_, new_n13750_, new_n13751_, new_n13752_, new_n13753_,
    new_n13754_, new_n13755_, new_n13756_, new_n13757_, new_n13758_,
    new_n13759_, new_n13760_, new_n13761_, new_n13762_, new_n13763_,
    new_n13764_, new_n13765_, new_n13766_, new_n13767_, new_n13768_,
    new_n13769_, new_n13770_, new_n13771_, new_n13772_, new_n13773_,
    new_n13774_, new_n13775_, new_n13776_, new_n13777_, new_n13778_,
    new_n13779_, new_n13780_, new_n13781_, new_n13782_, new_n13783_,
    new_n13784_, new_n13785_, new_n13786_, new_n13787_, new_n13788_,
    new_n13789_, new_n13790_, new_n13791_, new_n13792_, new_n13794_,
    new_n13795_, new_n13796_, new_n13797_, new_n13798_, new_n13799_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13815_, new_n13816_, new_n13817_,
    new_n13818_, new_n13819_, new_n13820_, new_n13822_, new_n13823_,
    new_n13824_, new_n13825_, new_n13826_, new_n13827_, new_n13829_,
    new_n13830_, new_n13831_, new_n13832_, new_n13833_, new_n13834_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13847_, new_n13849_, new_n13850_, new_n13851_, new_n13852_,
    new_n13853_, new_n13854_, new_n13856_, new_n13857_, new_n13858_,
    new_n13859_, new_n13860_, new_n13861_, new_n13863_, new_n13864_,
    new_n13865_, new_n13866_, new_n13867_, new_n13868_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13877_, new_n13878_, new_n13879_, new_n13880_, new_n13881_,
    new_n13882_, new_n13884_, new_n13885_, new_n13886_, new_n13887_,
    new_n13888_, new_n13889_, new_n13891_, new_n13892_, new_n13893_,
    new_n13894_, new_n13895_, new_n13896_, new_n13898_, new_n13899_,
    new_n13900_, new_n13901_, new_n13902_, new_n13903_, new_n13905_,
    new_n13906_, new_n13907_, new_n13908_, new_n13909_, new_n13910_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13919_, new_n13920_, new_n13921_, new_n13922_,
    new_n13923_, new_n13924_, new_n13926_, new_n13927_, new_n13928_,
    new_n13929_, new_n13930_, new_n13931_, new_n13933_, new_n13934_,
    new_n13935_, new_n13936_, new_n13937_, new_n13939_, new_n13940_,
    new_n13941_, new_n13942_, new_n13943_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13952_,
    new_n13953_, new_n13954_, new_n13955_, new_n13956_, new_n13957_,
    new_n13959_, new_n13960_, new_n13961_, new_n13962_, new_n13963_,
    new_n13965_, new_n13966_, new_n13967_, new_n13968_, new_n13969_,
    new_n13970_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13979_, new_n13980_, new_n13981_,
    new_n13982_, new_n13983_, new_n13984_, new_n13986_, new_n13987_,
    new_n13988_, new_n13989_, new_n13990_, new_n13991_, new_n13993_,
    new_n13994_, new_n13995_, new_n13996_, new_n13997_, new_n13998_,
    new_n14000_, new_n14001_, new_n14002_, new_n14003_, new_n14004_,
    new_n14005_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14012_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14020_, new_n14021_, new_n14022_,
    new_n14023_, new_n14024_, new_n14026_, new_n14027_, new_n14028_,
    new_n14029_, new_n14030_, new_n14032_, new_n14033_, new_n14034_,
    new_n14035_, new_n14036_, new_n14038_, new_n14039_, new_n14040_,
    new_n14041_, new_n14042_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14050_, new_n14051_, new_n14052_,
    new_n14053_, new_n14054_, new_n14056_, new_n14057_, new_n14058_,
    new_n14059_, new_n14060_, new_n14062_, new_n14063_, new_n14064_,
    new_n14065_, new_n14066_, new_n14068_, new_n14069_, new_n14070_,
    new_n14071_, new_n14072_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14080_, new_n14081_, new_n14082_,
    new_n14083_, new_n14084_, new_n14086_, new_n14087_, new_n14088_,
    new_n14089_, new_n14090_, new_n14092_, new_n14093_, new_n14094_,
    new_n14095_, new_n14096_, new_n14098_, new_n14099_, new_n14100_,
    new_n14101_, new_n14102_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14110_, new_n14111_, new_n14112_,
    new_n14113_, new_n14114_, new_n14116_, new_n14117_, new_n14118_,
    new_n14119_, new_n14120_, new_n14122_, new_n14123_, new_n14124_,
    new_n14125_, new_n14126_, new_n14128_, new_n14129_, new_n14130_,
    new_n14131_, new_n14132_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14140_, new_n14141_, new_n14142_,
    new_n14143_, new_n14144_, new_n14146_, new_n14147_, new_n14148_,
    new_n14149_, new_n14150_, new_n14151_, new_n14152_, new_n14153_,
    new_n14154_, new_n14155_, new_n14156_, new_n14157_, new_n14158_,
    new_n14159_, new_n14160_, new_n14161_, new_n14162_, new_n14163_,
    new_n14164_, new_n14166_, new_n14167_, new_n14168_, new_n14169_,
    new_n14170_, new_n14171_, new_n14172_, new_n14173_, new_n14174_,
    new_n14175_, new_n14176_, new_n14177_, new_n14178_, new_n14179_,
    new_n14180_, new_n14182_, new_n14183_, new_n14184_, new_n14185_,
    new_n14186_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14192_, new_n14193_, new_n14195_, new_n14196_, new_n14197_,
    new_n14198_, new_n14199_, new_n14201_, new_n14202_, new_n14203_,
    new_n14204_, new_n14205_, new_n14207_, new_n14208_, new_n14209_,
    new_n14210_, new_n14211_, new_n14212_, new_n14213_, new_n14214_,
    new_n14215_, new_n14216_, new_n14217_, new_n14218_, new_n14219_,
    new_n14220_, new_n14221_, new_n14222_, new_n14223_, new_n14224_,
    new_n14225_, new_n14226_, new_n14227_, new_n14228_, new_n14229_,
    new_n14230_, new_n14231_, new_n14232_, new_n14233_, new_n14234_,
    new_n14235_, new_n14236_, new_n14237_, new_n14238_, new_n14239_,
    new_n14240_, new_n14241_, new_n14242_, new_n14243_, new_n14244_,
    new_n14245_, new_n14246_, new_n14247_, new_n14248_, new_n14249_,
    new_n14250_, new_n14251_, new_n14252_, new_n14253_, new_n14254_,
    new_n14255_, new_n14256_, new_n14257_, new_n14258_, new_n14259_,
    new_n14260_, new_n14261_, new_n14262_, new_n14263_, new_n14264_,
    new_n14265_, new_n14266_, new_n14267_, new_n14268_, new_n14269_,
    new_n14270_, new_n14271_, new_n14272_, new_n14273_, new_n14274_,
    new_n14275_, new_n14276_, new_n14278_, new_n14279_, new_n14280_,
    new_n14281_, new_n14282_, new_n14283_, new_n14285_, new_n14286_,
    new_n14287_, new_n14288_, new_n14289_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14296_, new_n14297_,
    new_n14298_, new_n14300_, new_n14301_, new_n14302_, new_n14303_,
    new_n14304_, new_n14306_, new_n14307_, new_n14308_, new_n14309_,
    new_n14310_, new_n14312_, new_n14313_, new_n14314_, new_n14315_,
    new_n14316_, new_n14317_, new_n14319_, new_n14320_, new_n14321_,
    new_n14322_, new_n14323_, new_n14324_, new_n14326_, new_n14327_,
    new_n14328_, new_n14329_, new_n14330_, new_n14331_, new_n14333_,
    new_n14334_, new_n14335_, new_n14336_, new_n14337_, new_n14339_,
    new_n14340_, new_n14341_, new_n14342_, new_n14343_, new_n14345_,
    new_n14346_, new_n14347_, new_n14348_, new_n14349_, new_n14351_,
    new_n14352_, new_n14353_, new_n14354_, new_n14355_, new_n14357_,
    new_n14358_, new_n14359_, new_n14360_, new_n14361_, new_n14363_,
    new_n14364_, new_n14365_, new_n14366_, new_n14367_, new_n14368_,
    new_n14369_, new_n14371_, new_n14372_, new_n14373_, new_n14374_,
    new_n14375_, new_n14377_, new_n14378_, new_n14379_, new_n14380_,
    new_n14381_, new_n14383_, new_n14384_, new_n14385_, new_n14386_,
    new_n14388_, new_n14389_, new_n14390_, new_n14391_, new_n14392_,
    new_n14394_, new_n14395_, new_n14396_, new_n14397_, new_n14399_,
    new_n14400_, new_n14401_, new_n14402_, new_n14403_, new_n14405_,
    new_n14406_, new_n14407_, new_n14408_, new_n14409_, new_n14411_,
    new_n14412_, new_n14413_, new_n14414_, new_n14415_, new_n14417_,
    new_n14418_, new_n14419_, new_n14420_, new_n14421_, new_n14423_,
    new_n14424_, new_n14425_, new_n14426_, new_n14427_, new_n14428_,
    new_n14430_, new_n14431_, new_n14433_, new_n14434_, new_n14435_,
    new_n14436_, new_n14437_, new_n14438_, new_n14439_, new_n14440_,
    new_n14441_, new_n14442_, new_n14443_, new_n14444_, new_n14445_,
    new_n14446_, new_n14447_, new_n14448_, new_n14449_, new_n14450_,
    new_n14451_, new_n14452_, new_n14453_, new_n14454_, new_n14455_,
    new_n14456_, new_n14457_, new_n14458_, new_n14459_, new_n14460_,
    new_n14461_, new_n14462_, new_n14463_, new_n14464_, new_n14465_,
    new_n14466_, new_n14467_, new_n14468_, new_n14469_, new_n14470_,
    new_n14471_, new_n14472_, new_n14473_, new_n14474_, new_n14475_,
    new_n14476_, new_n14477_, new_n14478_, new_n14479_, new_n14480_,
    new_n14481_, new_n14482_, new_n14483_, new_n14484_, new_n14485_,
    new_n14486_, new_n14487_, new_n14488_, new_n14489_, new_n14490_,
    new_n14491_, new_n14492_, new_n14493_, new_n14494_, new_n14495_,
    new_n14496_, new_n14497_, new_n14498_, new_n14499_, new_n14500_,
    new_n14501_, new_n14502_, new_n14504_, new_n14505_, new_n14506_,
    new_n14507_, new_n14508_, new_n14509_, new_n14510_, new_n14511_,
    new_n14512_, new_n14513_, new_n14514_, new_n14515_, new_n14516_,
    new_n14517_, new_n14518_, new_n14519_, new_n14520_, new_n14521_,
    new_n14523_, new_n14524_, new_n14525_, new_n14526_, new_n14527_,
    new_n14528_, new_n14529_, new_n14530_, new_n14531_, new_n14532_,
    new_n14533_, new_n14534_, new_n14535_, new_n14536_, new_n14537_,
    new_n14538_, new_n14539_, new_n14540_, new_n14541_, new_n14542_,
    new_n14543_, new_n14544_, new_n14546_, new_n14547_, new_n14548_,
    new_n14549_, new_n14550_, new_n14551_, new_n14552_, new_n14553_,
    new_n14554_, new_n14555_, new_n14556_, new_n14557_, new_n14558_,
    new_n14559_, new_n14560_, new_n14561_, new_n14562_, new_n14563_,
    new_n14564_, new_n14565_, new_n14566_, new_n14567_, new_n14568_,
    new_n14569_, new_n14570_, new_n14571_, new_n14572_, new_n14573_,
    new_n14574_, new_n14575_, new_n14576_, new_n14577_, new_n14578_,
    new_n14579_, new_n14580_, new_n14581_, new_n14582_, new_n14583_,
    new_n14584_, new_n14585_, new_n14586_, new_n14587_, new_n14588_,
    new_n14589_, new_n14590_, new_n14591_, new_n14592_, new_n14593_,
    new_n14594_, new_n14595_, new_n14596_, new_n14597_, new_n14598_,
    new_n14599_, new_n14601_, new_n14602_, new_n14603_, new_n14604_,
    new_n14605_, new_n14606_, new_n14607_, new_n14608_, new_n14609_,
    new_n14610_, new_n14611_, new_n14612_, new_n14613_, new_n14614_,
    new_n14615_, new_n14616_, new_n14617_, new_n14618_, new_n14619_,
    new_n14620_, new_n14621_, new_n14622_, new_n14623_, new_n14624_,
    new_n14625_, new_n14627_, new_n14628_, new_n14629_, new_n14630_,
    new_n14631_, new_n14632_, new_n14633_, new_n14634_, new_n14635_,
    new_n14636_, new_n14637_, new_n14638_, new_n14639_, new_n14640_,
    new_n14641_, new_n14642_, new_n14643_, new_n14644_, new_n14645_,
    new_n14646_, new_n14647_, new_n14648_, new_n14649_, new_n14650_,
    new_n14651_, new_n14652_, new_n14653_, new_n14654_, new_n14656_,
    new_n14657_, new_n14658_, new_n14659_, new_n14660_, new_n14661_,
    new_n14662_, new_n14663_, new_n14664_, new_n14665_, new_n14666_,
    new_n14667_, new_n14668_, new_n14669_, new_n14670_, new_n14671_,
    new_n14672_, new_n14673_, new_n14674_, new_n14675_, new_n14676_,
    new_n14677_, new_n14678_, new_n14679_, new_n14680_, new_n14682_,
    new_n14683_, new_n14684_, new_n14685_, new_n14686_, new_n14687_,
    new_n14688_, new_n14689_, new_n14690_, new_n14691_, new_n14692_,
    new_n14693_, new_n14694_, new_n14695_, new_n14696_, new_n14697_,
    new_n14698_, new_n14700_, new_n14701_, new_n14702_, new_n14703_,
    new_n14704_, new_n14706_, new_n14707_, new_n14708_, new_n14709_,
    new_n14710_, new_n14711_, new_n14712_, new_n14713_, new_n14714_,
    new_n14715_, new_n14716_, new_n14717_, new_n14718_, new_n14719_,
    new_n14720_, new_n14721_, new_n14722_, new_n14723_, new_n14724_,
    new_n14725_, new_n14726_, new_n14727_, new_n14728_, new_n14729_,
    new_n14730_, new_n14731_, new_n14732_, new_n14734_, new_n14735_,
    new_n14736_, new_n14737_, new_n14738_, new_n14739_, new_n14740_,
    new_n14741_, new_n14742_, new_n14743_, new_n14744_, new_n14745_,
    new_n14746_, new_n14747_, new_n14748_, new_n14749_, new_n14751_,
    new_n14752_, new_n14753_, new_n14754_, new_n14755_, new_n14756_,
    new_n14757_, new_n14758_, new_n14759_, new_n14760_, new_n14761_,
    new_n14762_, new_n14763_, new_n14764_, new_n14765_, new_n14766_,
    new_n14768_, new_n14769_, new_n14770_, new_n14771_, new_n14772_,
    new_n14773_, new_n14774_, new_n14775_, new_n14776_, new_n14777_,
    new_n14778_, new_n14779_, new_n14780_, new_n14781_, new_n14782_,
    new_n14783_, new_n14784_, new_n14785_, new_n14786_, new_n14787_,
    new_n14788_, new_n14789_, new_n14790_, new_n14791_, new_n14792_,
    new_n14793_, new_n14794_, new_n14795_, new_n14796_, new_n14797_,
    new_n14798_, new_n14799_, new_n14801_, new_n14802_, new_n14803_,
    new_n14804_, new_n14805_, new_n14807_, new_n14808_, new_n14809_,
    new_n14810_, new_n14811_, new_n14812_, new_n14813_, new_n14814_,
    new_n14815_, new_n14816_, new_n14817_, new_n14818_, new_n14819_,
    new_n14820_, new_n14821_, new_n14822_, new_n14824_, new_n14825_,
    new_n14826_, new_n14827_, new_n14828_, new_n14829_, new_n14830_,
    new_n14831_, new_n14832_, new_n14833_, new_n14834_, new_n14835_,
    new_n14836_, new_n14837_, new_n14838_, new_n14839_, new_n14841_,
    new_n14842_, new_n14843_, new_n14844_, new_n14845_, new_n14847_,
    new_n14848_, new_n14849_, new_n14850_, new_n14851_, new_n14852_,
    new_n14853_, new_n14854_, new_n14855_, new_n14856_, new_n14857_,
    new_n14858_, new_n14859_, new_n14860_, new_n14861_, new_n14862_,
    new_n14864_, new_n14865_, new_n14866_, new_n14867_, new_n14868_,
    new_n14870_, new_n14871_, new_n14872_, new_n14873_, new_n14874_,
    new_n14875_, new_n14876_, new_n14878_, new_n14879_, new_n14880_,
    new_n14881_, new_n14882_, new_n14883_, new_n14884_, new_n14885_,
    new_n14886_, new_n14888_, new_n14889_, new_n14890_, new_n14891_,
    new_n14893_, new_n14894_, new_n14895_, new_n14896_, new_n14897_,
    new_n14898_, new_n14899_, new_n14900_, new_n14901_, new_n14902_,
    new_n14903_, new_n14904_, new_n14905_, new_n14907_, new_n14908_,
    new_n14909_, new_n14910_, new_n14911_, new_n14912_, new_n14913_,
    new_n14914_, new_n14915_, new_n14916_, new_n14917_, new_n14918_,
    new_n14919_, new_n14920_, new_n14921_, new_n14922_, new_n14923_,
    new_n14925_, new_n14926_, new_n14927_, new_n14928_, new_n14929_,
    new_n14931_, new_n14932_, new_n14933_, new_n14934_, new_n14935_,
    new_n14937_, new_n14938_, new_n14939_, new_n14940_, new_n14941_,
    new_n14943_, new_n14944_, new_n14945_, new_n14946_, new_n14947_,
    new_n14949_, new_n14950_, new_n14951_, new_n14952_, new_n14953_,
    new_n14955_, new_n14956_, new_n14957_, new_n14958_, new_n14959_,
    new_n14961_, new_n14962_, new_n14963_, new_n14964_, new_n14965_,
    new_n14967_, new_n14968_, new_n14969_, new_n14970_, new_n14971_,
    new_n14972_, new_n14973_, new_n14974_, new_n14975_, new_n14976_,
    new_n14977_, new_n14979_, new_n14980_, new_n14981_, new_n14982_,
    new_n14983_, new_n14984_, new_n14985_, new_n14986_, new_n14987_,
    new_n14988_, new_n14989_, new_n14990_, new_n14991_, new_n14992_,
    new_n14993_, new_n14994_, new_n14995_, new_n14997_, new_n14998_,
    new_n14999_, new_n15000_, new_n15001_, new_n15002_, new_n15003_,
    new_n15004_, new_n15005_, new_n15006_, new_n15008_, new_n15009_,
    new_n15010_, new_n15011_, new_n15012_, new_n15013_, new_n15014_,
    new_n15015_, new_n15016_, new_n15017_, new_n15019_, new_n15020_,
    new_n15021_, new_n15022_, new_n15023_, new_n15024_, new_n15025_,
    new_n15026_, new_n15027_, new_n15028_, new_n15030_, new_n15031_,
    new_n15032_, new_n15033_, new_n15034_, new_n15035_, new_n15036_,
    new_n15037_, new_n15038_, new_n15039_, new_n15040_, new_n15041_,
    new_n15042_, new_n15043_, new_n15044_, new_n15045_, new_n15046_,
    new_n15047_, new_n15048_, new_n15050_, new_n15051_, new_n15052_,
    new_n15053_, new_n15054_, new_n15055_, new_n15056_, new_n15057_,
    new_n15058_, new_n15059_, new_n15060_, new_n15061_, new_n15062_,
    new_n15064_, new_n15065_, new_n15066_, new_n15067_, new_n15068_,
    new_n15069_, new_n15070_, new_n15071_, new_n15072_, new_n15073_,
    new_n15075_, new_n15076_, new_n15077_, new_n15078_, new_n15079_,
    new_n15080_, new_n15081_, new_n15082_, new_n15083_, new_n15084_,
    new_n15086_, new_n15087_, new_n15088_, new_n15089_, new_n15090_,
    new_n15091_, new_n15092_, new_n15093_, new_n15094_, new_n15095_,
    new_n15096_, new_n15097_, new_n15098_, new_n15100_, new_n15101_,
    new_n15102_, new_n15103_, new_n15104_, new_n15105_, new_n15106_,
    new_n15107_, new_n15108_, new_n15109_, new_n15110_, new_n15111_,
    new_n15112_, new_n15114_, new_n15115_, new_n15116_, new_n15117_,
    new_n15118_, new_n15119_, new_n15120_, new_n15121_, new_n15122_,
    new_n15123_, new_n15124_, new_n15125_, new_n15126_, new_n15128_,
    new_n15129_, new_n15130_, new_n15131_, new_n15132_, new_n15133_,
    new_n15134_, new_n15135_, new_n15136_, new_n15137_, new_n15139_,
    new_n15140_, new_n15141_, new_n15142_, new_n15143_, new_n15144_,
    new_n15145_, new_n15146_, new_n15147_, new_n15148_, new_n15149_,
    new_n15150_, new_n15151_, new_n15153_, new_n15154_, new_n15155_,
    new_n15156_, new_n15157_, new_n15158_, new_n15159_, new_n15160_,
    new_n15161_, new_n15162_, new_n15163_, new_n15164_, new_n15165_,
    new_n15167_, new_n15168_, new_n15169_, new_n15170_, new_n15171_,
    new_n15172_, new_n15173_, new_n15174_, new_n15175_, new_n15176_,
    new_n15178_, new_n15179_, new_n15180_, new_n15181_, new_n15182_,
    new_n15183_, new_n15184_, new_n15185_, new_n15186_, new_n15187_,
    new_n15189_, new_n15190_, new_n15191_, new_n15192_, new_n15193_,
    new_n15194_, new_n15195_, new_n15196_, new_n15197_, new_n15198_,
    new_n15200_, new_n15201_, new_n15202_, new_n15203_, new_n15204_,
    new_n15205_, new_n15206_, new_n15207_, new_n15208_, new_n15209_,
    new_n15211_, new_n15212_, new_n15213_, new_n15214_, new_n15215_,
    new_n15216_, new_n15217_, new_n15218_, new_n15219_, new_n15220_,
    new_n15222_, new_n15223_, new_n15224_, new_n15225_, new_n15226_,
    new_n15227_, new_n15228_, new_n15229_, new_n15230_, new_n15231_,
    new_n15233_, new_n15234_, new_n15235_, new_n15236_, new_n15237_,
    new_n15238_, new_n15239_, new_n15240_, new_n15241_, new_n15242_,
    new_n15243_, new_n15244_, new_n15245_, new_n15247_, new_n15248_,
    new_n15249_, new_n15250_, new_n15252_, new_n15253_, new_n15254_,
    new_n15255_, new_n15256_, new_n15257_, new_n15258_, new_n15259_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15266_, new_n15268_, new_n15269_, new_n15270_,
    new_n15271_, new_n15272_, new_n15273_, new_n15274_, new_n15275_,
    new_n15276_, new_n15277_, new_n15279_, new_n15281_, new_n15282_,
    new_n15283_, new_n15284_, new_n15285_, new_n15286_, new_n15288_,
    new_n15289_, new_n15290_, new_n15291_, new_n15292_, new_n15293_,
    new_n15294_, new_n15295_, new_n15296_, new_n15297_, new_n15299_,
    new_n15300_, new_n15302_, new_n15303_, new_n15305_, new_n15306_,
    new_n15308_, new_n15309_, new_n15311_, new_n15312_, new_n15314_,
    new_n15315_, new_n15317_, new_n15318_, new_n15320_, new_n15321_,
    new_n15323_, new_n15324_, new_n15326_, new_n15327_, new_n15328_,
    new_n15329_, new_n15330_, new_n15331_, new_n15332_, new_n15333_,
    new_n15334_, new_n15335_, new_n15336_, new_n15337_, new_n15338_,
    new_n15339_, new_n15340_, new_n15341_, new_n15342_, new_n15343_,
    new_n15344_, new_n15345_, new_n15346_, new_n15347_, new_n15348_,
    new_n15349_, new_n15350_, new_n15351_, new_n15353_, new_n15354_,
    new_n15355_, new_n15356_, new_n15357_, new_n15358_, new_n15360_,
    new_n15361_, new_n15362_, new_n15363_, new_n15364_, new_n15365_,
    new_n15367_, new_n15368_, new_n15369_, new_n15370_, new_n15371_,
    new_n15372_, new_n15373_, new_n15375_, new_n15376_, new_n15378_,
    new_n15379_, new_n15381_, new_n15382_, new_n15384_, new_n15385_,
    new_n15387_, new_n15388_, new_n15390_, new_n15391_, new_n15393_,
    new_n15394_, new_n15396_, new_n15397_, new_n15398_, new_n15399_,
    new_n15400_, new_n15401_, new_n15402_, new_n15404_, new_n15405_,
    new_n15406_, new_n15407_, new_n15408_, new_n15409_, new_n15411_,
    new_n15412_, new_n15413_, new_n15415_, new_n15416_, new_n15417_,
    new_n15418_, new_n15419_, new_n15421_, new_n15422_, new_n15424_,
    new_n15425_, new_n15426_, new_n15427_, new_n15429_, new_n15430_,
    new_n15431_, new_n15433_, new_n15434_, new_n15436_, new_n15437_,
    new_n15438_, new_n15440_, new_n15441_, new_n15442_, new_n15444_,
    new_n15445_, new_n15447_, new_n15448_, new_n15450_, new_n15451_,
    new_n15453_, new_n15454_, new_n15456_, new_n15457_, new_n15459_,
    new_n15460_, new_n15462_, new_n15463_, new_n15465_, new_n15466_,
    new_n15468_, new_n15469_, new_n15471_, new_n15472_, new_n15474_,
    new_n15475_, new_n15477_, new_n15478_, new_n15479_, new_n15481_,
    new_n15482_, new_n15484_, new_n15486_, new_n15487_, new_n15489_,
    new_n15490_, new_n15492_, new_n15493_, new_n15495_, new_n15496_,
    new_n15498_, new_n15499_, new_n15501_, new_n15502_, new_n15504_,
    new_n15505_, new_n15507_, new_n15508_, new_n15509_, new_n15511_,
    new_n15512_, new_n15514_, new_n15515_, new_n15517_, new_n15518_,
    new_n15520_, new_n15521_, new_n15523_, new_n15524_, new_n15526_,
    new_n15527_, new_n15529_, new_n15530_, new_n15532_, new_n15533_,
    new_n15535_, new_n15536_, new_n15538_, new_n15539_, new_n15541_,
    new_n15542_, new_n15544_, new_n15545_, new_n15547_, new_n15548_,
    new_n15550_, new_n15551_, new_n15553_, new_n15554_, new_n15556_,
    new_n15557_, new_n15559_, new_n15560_, new_n15562_, new_n15563_,
    new_n15565_, new_n15566_, new_n15568_, new_n15569_, new_n15571_,
    new_n15572_, new_n15574_, new_n15575_, new_n15577_, new_n15578_,
    new_n15580_, new_n15581_, new_n15583_, new_n15584_, new_n15586_,
    new_n15587_, new_n15589_, new_n15590_, new_n15592_, new_n15593_,
    new_n15595_, new_n15596_, new_n15598_, new_n15599_, new_n15601_,
    new_n15602_, new_n15604_, new_n15605_, new_n15607_, new_n15608_,
    new_n15610_, new_n15611_, new_n15613_, new_n15614_, new_n15616_,
    new_n15617_, new_n15619_, new_n15620_, new_n15622_, new_n15623_,
    new_n15625_, new_n15626_, new_n15628_, new_n15629_, new_n15631_,
    new_n15632_, new_n15634_, new_n15635_, new_n15637_, new_n15638_,
    new_n15640_, new_n15641_, new_n15643_, new_n15644_, new_n15646_,
    new_n15647_, new_n15649_, new_n15650_, new_n15652_, new_n15653_,
    new_n15655_, new_n15656_, new_n15658_, new_n15659_, new_n15661_,
    new_n15662_, new_n15664_, new_n15665_, new_n15667_, new_n15668_,
    new_n15670_, new_n15671_, new_n15673_, new_n15674_, new_n15676_,
    new_n15677_, new_n15679_, new_n15680_, new_n15682_, new_n15683_,
    new_n15685_, new_n15686_, new_n15688_, new_n15689_, new_n15691_,
    new_n15692_, new_n15694_, new_n15695_, new_n15697_, new_n15698_,
    new_n15700_, new_n15701_, new_n15703_, new_n15704_, new_n15706_,
    new_n15707_, new_n15709_, new_n15710_, new_n15712_, new_n15713_,
    new_n15715_, new_n15716_, new_n15718_, new_n15719_, new_n15721_,
    new_n15722_, new_n15724_, new_n15725_, new_n15727_, new_n15728_,
    new_n15730_, new_n15731_, new_n15733_, new_n15734_, new_n15736_,
    new_n15737_, new_n15739_, new_n15740_, new_n15742_, new_n15743_,
    new_n15745_, new_n15746_, new_n15748_, new_n15749_, new_n15751_,
    new_n15752_, new_n15754_, new_n15755_, new_n15757_, new_n15758_,
    new_n15760_, new_n15761_, new_n15763_, new_n15764_, new_n15766_,
    new_n15767_, new_n15769_, new_n15770_, new_n15772_, new_n15773_,
    new_n15775_, new_n15776_, new_n15778_, new_n15779_, new_n15781_,
    new_n15782_, new_n15784_, new_n15785_, new_n15787_, new_n15788_,
    new_n15790_, new_n15791_, new_n15793_, new_n15794_, new_n15796_,
    new_n15797_, new_n15799_, new_n15800_, new_n15802_, new_n15803_,
    new_n15805_, new_n15806_, new_n15808_, new_n15809_, new_n15811_,
    new_n15812_, new_n15814_, new_n15815_, new_n15817_, new_n15818_,
    new_n15820_, new_n15821_, new_n15823_, new_n15824_, new_n15826_,
    new_n15827_, new_n15829_, new_n15830_, new_n15832_, new_n15833_,
    new_n15835_, new_n15836_, new_n15838_, new_n15839_, new_n15841_,
    new_n15842_, new_n15844_, new_n15845_, new_n15847_, new_n15848_,
    new_n15850_, new_n15851_, new_n15853_, new_n15854_, new_n15856_,
    new_n15857_, new_n15859_, new_n15860_, new_n15861_, new_n15862_,
    new_n15863_, new_n15864_, new_n15865_, new_n15866_, new_n15867_,
    new_n15868_, new_n15869_, new_n15870_, new_n15871_, new_n15872_,
    new_n15873_, new_n15874_, new_n15875_, new_n15876_, new_n15877_,
    new_n15878_, new_n15879_, new_n15880_, new_n15881_, new_n15882_,
    new_n15883_, new_n15884_, new_n15885_, new_n15886_, new_n15887_,
    new_n15888_, new_n15889_, new_n15890_, new_n15891_, new_n15892_,
    new_n15893_, new_n15894_, new_n15895_, new_n15896_, new_n15897_,
    new_n15898_, new_n15899_, new_n15900_, new_n15901_, new_n15902_,
    new_n15903_, new_n15904_, new_n15905_, new_n15906_, new_n15907_,
    new_n15908_, new_n15909_, new_n15910_, new_n15912_, new_n15913_,
    new_n15915_, new_n15916_, new_n15918_, new_n15919_, new_n15921_,
    new_n15922_, new_n15924_, new_n15925_, new_n15927_, new_n15928_,
    new_n15930_, new_n15931_, new_n15933_, new_n15934_, new_n15935_,
    new_n15936_, new_n15937_, new_n15939_, new_n15940_, new_n15941_,
    new_n15942_, new_n15943_, new_n15945_, new_n15946_, new_n15947_,
    new_n15948_, new_n15949_, new_n15950_, new_n15951_, new_n15952_,
    new_n15953_, new_n15954_, new_n15955_, new_n15956_, new_n15957_,
    new_n15958_, new_n15959_, new_n15960_, new_n15961_, new_n15962_,
    new_n15963_, new_n15964_, new_n15965_, new_n15966_, new_n15967_,
    new_n15968_, new_n15969_, new_n15970_, new_n15971_, new_n15973_,
    new_n15974_, new_n15975_, new_n15977_, new_n15978_, new_n15979_,
    new_n15980_, new_n15981_, new_n15983_, new_n15984_, new_n15985_,
    new_n15986_, new_n15987_, new_n15989_, new_n15990_, new_n15991_,
    new_n15992_, new_n15993_, new_n15995_, new_n15996_, new_n15997_,
    new_n15998_, new_n15999_, new_n16001_, new_n16002_, new_n16003_,
    new_n16004_, new_n16005_, new_n16007_, new_n16008_, new_n16009_,
    new_n16010_, new_n16011_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16019_, new_n16020_, new_n16021_,
    new_n16022_, new_n16023_, new_n16024_, new_n16025_, new_n16026_,
    new_n16027_, new_n16028_, new_n16029_, new_n16030_, new_n16031_,
    new_n16032_, new_n16033_, new_n16034_, new_n16035_, new_n16036_,
    new_n16037_, new_n16038_, new_n16039_, new_n16040_, new_n16041_,
    new_n16042_, new_n16045_, new_n16046_, new_n16048_, new_n16049_,
    new_n16051_, new_n16052_, new_n16054_, new_n16055_, new_n16057_,
    new_n16058_, new_n16060_, new_n16061_, new_n16063_, new_n16064_,
    new_n16066_, new_n16067_, new_n16069_, new_n16070_, new_n16072_,
    new_n16073_, new_n16075_, new_n16076_, new_n16078_, new_n16079_,
    new_n16081_, new_n16082_, new_n16084_, new_n16085_, new_n16087_,
    new_n16088_, new_n16090_, new_n16091_, new_n16093_, new_n16094_,
    new_n16096_, new_n16097_, new_n16099_, new_n16100_, new_n16102_,
    new_n16103_, new_n16105_, new_n16106_, new_n16108_, new_n16109_,
    new_n16111_, new_n16112_, new_n16114_, new_n16115_, new_n16117_,
    new_n16118_, new_n16120_, new_n16121_, new_n16123_, new_n16124_,
    new_n16126_, new_n16127_, new_n16129_, new_n16130_, new_n16132_,
    new_n16133_, new_n16135_, new_n16136_, new_n16138_, new_n16139_,
    new_n16141_, new_n16142_, new_n16144_, new_n16145_, new_n16147_,
    new_n16148_, new_n16150_, new_n16151_, new_n16153_, new_n16154_,
    new_n16156_, new_n16157_, new_n16159_, new_n16160_, new_n16162_,
    new_n16163_, new_n16165_, new_n16166_, new_n16168_, new_n16169_,
    new_n16171_, new_n16172_, new_n16174_, new_n16175_, new_n16177_,
    new_n16178_, new_n16180_, new_n16181_, new_n16183_, new_n16184_,
    new_n16186_, new_n16187_, new_n16189_, new_n16190_, new_n16192_,
    new_n16193_, new_n16195_, new_n16196_, new_n16198_, new_n16199_,
    new_n16201_, new_n16202_, new_n16204_, new_n16205_, new_n16207_,
    new_n16208_, new_n16210_, new_n16211_, new_n16213_, new_n16214_,
    new_n16216_, new_n16217_, new_n16219_, new_n16220_, new_n16222_,
    new_n16223_, new_n16225_, new_n16226_, new_n16228_, new_n16229_,
    new_n16231_, new_n16232_, new_n16234_, new_n16235_, new_n16237_,
    new_n16238_, new_n16240_, new_n16241_, new_n16243_, new_n16244_,
    new_n16246_, new_n16247_, new_n16249_, new_n16250_, new_n16252_,
    new_n16253_, new_n16255_, new_n16256_, new_n16258_, new_n16259_,
    new_n16261_, new_n16262_, new_n16264_, new_n16265_, new_n16267_,
    new_n16268_, new_n16270_, new_n16271_, new_n16273_, new_n16274_,
    new_n16276_, new_n16277_, new_n16279_, new_n16280_, new_n16282_,
    new_n16283_, new_n16285_, new_n16286_, new_n16288_, new_n16289_,
    new_n16291_, new_n16292_, new_n16294_, new_n16295_, new_n16297_,
    new_n16298_, new_n16300_, new_n16301_, new_n16304_, new_n16305_,
    new_n16306_, new_n16307_, new_n16308_, new_n16309_, new_n16310_,
    new_n16312_, new_n16313_, new_n16315_, new_n16316_, new_n16318_,
    new_n16319_, new_n16321_, new_n16322_, new_n16324_, new_n16325_,
    new_n16327_, new_n16328_, new_n16330_, new_n16331_, new_n16333_,
    new_n16334_, new_n16336_, new_n16337_, new_n16339_, new_n16340_,
    new_n16342_, new_n16343_, new_n16345_, new_n16346_, new_n16348_,
    new_n16349_, new_n16351_, new_n16352_, new_n16354_, new_n16355_,
    new_n16357_, new_n16358_, new_n16360_, new_n16361_, new_n16363_,
    new_n16364_, new_n16366_, new_n16367_, new_n16369_, new_n16370_,
    new_n16371_, new_n16372_, new_n16374_, new_n16375_, new_n16376_,
    new_n16377_, new_n16378_, new_n16379_, new_n16380_, new_n16381_,
    new_n16382_, new_n16383_, new_n16384_, new_n16385_, new_n16386_,
    new_n16387_, new_n16388_, new_n16389_, new_n16391_, new_n16392_,
    new_n16393_, new_n16395_, new_n16396_, new_n16397_, new_n16399_,
    new_n16400_, new_n16401_, new_n16403_, new_n16404_, new_n16405_,
    new_n16406_, new_n16407_, new_n16408_, new_n16409_, new_n16410_,
    new_n16411_, new_n16412_, new_n16413_, new_n16414_, new_n16415_,
    new_n16416_, new_n16417_, new_n16418_, new_n16419_, new_n16420_,
    new_n16421_, new_n16422_, new_n16423_, new_n16424_, new_n16425_,
    new_n16426_, new_n16427_, new_n16428_, new_n16429_, new_n16430_,
    new_n16431_, new_n16432_, new_n16433_, new_n16434_, new_n16435_,
    new_n16436_, new_n16437_, new_n16438_, new_n16439_, new_n16440_,
    new_n16441_, new_n16442_, new_n16443_, new_n16444_, new_n16445_,
    new_n16446_, new_n16447_, new_n16448_, new_n16449_, new_n16450_,
    new_n16451_, new_n16452_, new_n16453_, new_n16454_, new_n16455_,
    new_n16456_, new_n16457_, new_n16458_, new_n16459_, new_n16460_,
    new_n16461_, new_n16462_, new_n16463_, new_n16464_, new_n16465_,
    new_n16466_, new_n16467_, new_n16468_, new_n16469_, new_n16470_,
    new_n16471_, new_n16472_, new_n16473_, new_n16474_, new_n16475_,
    new_n16476_, new_n16477_, new_n16478_, new_n16479_, new_n16480_,
    new_n16481_, new_n16482_, new_n16483_, new_n16484_, new_n16485_,
    new_n16486_, new_n16487_, new_n16488_, new_n16489_, new_n16490_,
    new_n16491_, new_n16492_, new_n16493_, new_n16494_, new_n16495_,
    new_n16496_, new_n16497_, new_n16498_, new_n16499_, new_n16500_,
    new_n16501_, new_n16502_, new_n16503_, new_n16504_, new_n16505_,
    new_n16506_, new_n16507_, new_n16508_, new_n16509_, new_n16510_,
    new_n16511_, new_n16512_, new_n16513_, new_n16514_, new_n16515_,
    new_n16516_, new_n16517_, new_n16518_, new_n16519_, new_n16520_,
    new_n16521_, new_n16522_, new_n16523_, new_n16524_, new_n16525_,
    new_n16526_, new_n16527_, new_n16528_, new_n16529_, new_n16530_,
    new_n16531_, new_n16532_, new_n16533_, new_n16534_, new_n16535_,
    new_n16536_, new_n16537_, new_n16538_, new_n16539_, new_n16540_,
    new_n16541_, new_n16542_, new_n16543_, new_n16544_, new_n16545_,
    new_n16546_, new_n16547_, new_n16548_, new_n16549_, new_n16550_,
    new_n16551_, new_n16552_, new_n16553_, new_n16554_, new_n16555_,
    new_n16556_, new_n16557_, new_n16558_, new_n16559_, new_n16560_,
    new_n16561_, new_n16562_, new_n16563_, new_n16564_, new_n16565_,
    new_n16566_, new_n16567_, new_n16568_, new_n16569_, new_n16570_,
    new_n16571_, new_n16572_, new_n16573_, new_n16574_, new_n16575_,
    new_n16576_, new_n16577_, new_n16578_, new_n16579_, new_n16580_,
    new_n16581_, new_n16582_, new_n16583_, new_n16584_, new_n16585_,
    new_n16586_, new_n16587_, new_n16588_, new_n16589_, new_n16590_,
    new_n16591_, new_n16592_, new_n16593_, new_n16594_, new_n16595_,
    new_n16596_, new_n16597_, new_n16598_, new_n16599_, new_n16600_,
    new_n16601_, new_n16602_, new_n16603_, new_n16604_, new_n16605_,
    new_n16606_, new_n16607_, new_n16608_, new_n16609_, new_n16610_,
    new_n16611_, new_n16612_, new_n16613_, new_n16614_, new_n16615_,
    new_n16616_, new_n16617_, new_n16618_, new_n16619_, new_n16620_,
    new_n16621_, new_n16622_, new_n16623_, new_n16624_, new_n16625_,
    new_n16626_, new_n16627_, new_n16628_, new_n16629_, new_n16630_,
    new_n16631_, new_n16632_, new_n16633_, new_n16634_, new_n16635_,
    new_n16636_, new_n16637_, new_n16638_, new_n16639_, new_n16640_,
    new_n16641_, new_n16642_, new_n16643_, new_n16644_, new_n16645_,
    new_n16646_, new_n16647_, new_n16648_, new_n16649_, new_n16650_,
    new_n16651_, new_n16652_, new_n16653_, new_n16654_, new_n16655_,
    new_n16656_, new_n16657_, new_n16658_, new_n16659_, new_n16660_,
    new_n16661_, new_n16662_, new_n16663_, new_n16664_, new_n16665_,
    new_n16666_, new_n16667_, new_n16668_, new_n16669_, new_n16670_,
    new_n16671_, new_n16672_, new_n16673_, new_n16674_, new_n16675_,
    new_n16676_, new_n16677_, new_n16678_, new_n16679_, new_n16680_,
    new_n16681_, new_n16682_, new_n16683_, new_n16684_, new_n16685_,
    new_n16686_, new_n16687_, new_n16688_, new_n16689_, new_n16690_,
    new_n16691_, new_n16692_, new_n16693_, new_n16694_, new_n16695_,
    new_n16696_, new_n16697_, new_n16698_, new_n16699_, new_n16700_,
    new_n16701_, new_n16702_, new_n16703_, new_n16704_, new_n16705_,
    new_n16706_, new_n16707_, new_n16708_, new_n16709_, new_n16710_,
    new_n16711_, new_n16712_, new_n16713_, new_n16714_, new_n16715_,
    new_n16716_, new_n16717_, new_n16718_, new_n16719_, new_n16720_,
    new_n16721_, new_n16722_, new_n16723_, new_n16724_, new_n16725_,
    new_n16726_, new_n16727_, new_n16728_, new_n16729_, new_n16730_,
    new_n16731_, new_n16732_, new_n16733_, new_n16735_, new_n16736_,
    new_n16737_, new_n16738_, new_n16739_, new_n16741_, new_n16742_,
    new_n16743_, new_n16744_, new_n16745_, new_n16746_, new_n16747_,
    new_n16748_, new_n16750_, new_n16751_, new_n16752_, new_n16753_,
    new_n16754_, new_n16755_, new_n16756_, new_n16757_, new_n16759_,
    new_n16760_, new_n16761_, new_n16762_, new_n16763_, new_n16764_,
    new_n16767_, new_n16768_, new_n16769_, new_n16770_, new_n16771_,
    new_n16772_, new_n16774_, new_n16775_, new_n16776_, new_n16777_,
    new_n16778_, new_n16779_, new_n16780_, new_n16781_, new_n16783_,
    new_n16784_, new_n16785_, new_n16786_, new_n16787_, new_n16789_,
    new_n16790_, new_n16791_, new_n16792_, new_n16793_, new_n16794_,
    new_n16796_, new_n16797_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16805_, new_n16806_, new_n16807_,
    new_n16808_, new_n16809_, new_n16810_, new_n16812_, new_n16813_,
    new_n16814_, new_n16815_, new_n16816_, new_n16817_, new_n16818_,
    new_n16820_, new_n16821_, new_n16822_, new_n16824_, new_n16825_,
    new_n16826_, new_n16827_, new_n16828_, new_n16830_, new_n16831_,
    new_n16832_, new_n16834_, new_n16835_, new_n16836_, new_n16838_,
    new_n16839_, new_n16840_, new_n16842_, new_n16843_, new_n16844_,
    new_n16846_, new_n16847_, new_n16848_, new_n16850_, new_n16851_,
    new_n16852_, new_n16854_, new_n16855_, new_n16856_, new_n16858_,
    new_n16859_, new_n16860_, new_n16861_, new_n16863_, new_n16864_,
    new_n16865_, new_n16866_, new_n16867_, new_n16869_, new_n16870_,
    new_n16871_, new_n16872_, new_n16874_, new_n16875_, new_n16876_,
    new_n16877_, new_n16878_, new_n16880_, new_n16881_, new_n16882_,
    new_n16884_, new_n16885_, new_n16886_, new_n16888_, new_n16889_,
    new_n16890_, new_n16892_, new_n16893_, new_n16894_, new_n16896_,
    new_n16897_, new_n16898_, new_n16900_, new_n16901_, new_n16902_,
    new_n16904_, new_n16905_, new_n16906_, new_n16907_, new_n16908_,
    new_n16910_, new_n16911_, new_n16912_, new_n16913_, new_n16915_,
    new_n16916_, new_n16917_, new_n16919_, new_n16920_, new_n16921_,
    new_n16923_, new_n16924_, new_n16925_, new_n16927_, new_n16928_,
    new_n16929_, new_n16931_, new_n16932_, new_n16933_, new_n16935_,
    new_n16936_, new_n16937_, new_n16939_, new_n16940_, new_n16941_,
    new_n16943_, new_n16944_, new_n16945_, new_n16947_, new_n16948_,
    new_n16949_, new_n16951_, new_n16952_, new_n16953_, new_n16955_,
    new_n16956_, new_n16957_, new_n16959_, new_n16960_, new_n16961_,
    new_n16963_, new_n16964_, new_n16965_, new_n16967_, new_n16968_,
    new_n16969_, new_n16971_, new_n16972_, new_n16973_, new_n16975_,
    new_n16976_, new_n16977_, new_n16979_, new_n16980_, new_n16981_,
    new_n16983_, new_n16984_, new_n16985_, new_n16987_, new_n16988_,
    new_n16989_, new_n16991_, new_n16992_, new_n16993_, new_n16995_,
    new_n16996_, new_n16997_, new_n16999_, new_n17000_, new_n17001_,
    new_n17003_, new_n17004_, new_n17005_, new_n17007_, new_n17008_,
    new_n17009_, new_n17011_, new_n17012_, new_n17013_, new_n17015_,
    new_n17016_, new_n17017_, new_n17019_, new_n17020_, new_n17021_,
    new_n17023_, new_n17024_, new_n17025_, new_n17027_, new_n17028_,
    new_n17029_, new_n17031_, new_n17032_, new_n17033_, new_n17035_,
    new_n17036_, new_n17037_, new_n17039_, new_n17040_, new_n17041_,
    new_n17043_, new_n17044_, new_n17045_, new_n17047_, new_n17048_,
    new_n17049_, new_n17051_, new_n17052_, new_n17053_, new_n17054_,
    new_n17055_, new_n17056_, new_n17057_, new_n17058_, new_n17059_,
    new_n17060_, new_n17061_, new_n17062_, new_n17064_, new_n17065_,
    new_n17066_, new_n17068_, new_n17069_, new_n17070_, new_n17072_,
    new_n17073_, new_n17074_, new_n17076_, new_n17077_, new_n17078_,
    new_n17079_, new_n17080_, new_n17081_, new_n17082_, new_n17083_,
    new_n17084_, new_n17085_, new_n17086_, new_n17087_, new_n17088_,
    new_n17089_, new_n17090_, new_n17091_, new_n17092_, new_n17093_,
    new_n17094_, new_n17095_, new_n17096_, new_n17097_, new_n17098_,
    new_n17099_, new_n17100_, new_n17101_, new_n17102_, new_n17103_,
    new_n17104_, new_n17105_, new_n17106_, new_n17107_, new_n17108_,
    new_n17109_, new_n17110_, new_n17111_, new_n17112_, new_n17113_,
    new_n17114_, new_n17115_, new_n17116_, new_n17117_, new_n17118_,
    new_n17120_, new_n17121_, new_n17122_, new_n17123_, new_n17124_,
    new_n17125_, new_n17126_, new_n17127_, new_n17128_, new_n17129_,
    new_n17130_, new_n17131_, new_n17132_, new_n17133_, new_n17134_,
    new_n17135_, new_n17136_, new_n17137_, new_n17138_, new_n17139_,
    new_n17140_, new_n17142_, new_n17143_, new_n17144_, new_n17146_,
    new_n17147_, new_n17148_, new_n17149_, new_n17150_, new_n17151_,
    new_n17152_, new_n17153_, new_n17154_, new_n17155_, new_n17156_,
    new_n17157_, new_n17158_, new_n17159_, new_n17160_, new_n17161_,
    new_n17162_, new_n17163_, new_n17164_, new_n17165_, new_n17166_,
    new_n17168_, new_n17169_, new_n17170_, new_n17171_, new_n17172_,
    new_n17173_, new_n17174_, new_n17175_, new_n17176_, new_n17177_,
    new_n17178_, new_n17179_, new_n17180_, new_n17181_, new_n17182_,
    new_n17183_, new_n17184_, new_n17185_, new_n17186_, new_n17187_,
    new_n17188_, new_n17190_, new_n17191_, new_n17192_, new_n17193_,
    new_n17194_, new_n17195_, new_n17196_, new_n17197_, new_n17198_,
    new_n17199_, new_n17200_, new_n17201_, new_n17202_, new_n17203_,
    new_n17204_, new_n17205_, new_n17206_, new_n17207_, new_n17208_,
    new_n17209_, new_n17210_, new_n17212_, new_n17213_, new_n17214_,
    new_n17216_, new_n17217_, new_n17218_, new_n17219_, new_n17220_,
    new_n17221_, new_n17222_, new_n17223_, new_n17224_, new_n17225_,
    new_n17226_, new_n17227_, new_n17228_, new_n17229_, new_n17230_,
    new_n17231_, new_n17232_, new_n17234_, new_n17235_, new_n17236_,
    new_n17237_, new_n17238_, new_n17239_, new_n17240_, new_n17241_,
    new_n17242_, new_n17243_, new_n17244_, new_n17245_, new_n17246_,
    new_n17247_, new_n17248_, new_n17249_, new_n17250_, new_n17252_,
    new_n17253_, new_n17254_, new_n17255_, new_n17256_, new_n17257_,
    new_n17258_, new_n17259_, new_n17260_, new_n17261_, new_n17262_,
    new_n17263_, new_n17264_, new_n17265_, new_n17266_, new_n17267_,
    new_n17268_, new_n17269_, new_n17270_, new_n17271_, new_n17272_,
    new_n17274_, new_n17275_, new_n17276_, new_n17277_, new_n17278_,
    new_n17279_, new_n17280_, new_n17281_, new_n17282_, new_n17283_,
    new_n17284_, new_n17285_, new_n17286_, new_n17287_, new_n17288_,
    new_n17289_, new_n17290_, new_n17291_, new_n17292_, new_n17293_,
    new_n17294_, new_n17296_, new_n17297_, new_n17298_, new_n17299_,
    new_n17300_, new_n17301_, new_n17302_, new_n17303_, new_n17304_,
    new_n17305_, new_n17306_, new_n17307_, new_n17308_, new_n17309_,
    new_n17310_, new_n17311_, new_n17312_, new_n17313_, new_n17314_,
    new_n17315_, new_n17316_, new_n17318_, new_n17319_, new_n17320_,
    new_n17321_, new_n17322_, new_n17323_, new_n17324_, new_n17325_,
    new_n17326_, new_n17327_, new_n17328_, new_n17329_, new_n17330_,
    new_n17331_, new_n17332_, new_n17333_, new_n17334_, new_n17335_,
    new_n17336_, new_n17337_, new_n17338_, new_n17340_, new_n17341_,
    new_n17342_, new_n17343_, new_n17344_, new_n17345_, new_n17346_,
    new_n17347_, new_n17348_, new_n17349_, new_n17350_, new_n17351_,
    new_n17352_, new_n17353_, new_n17354_, new_n17355_, new_n17356_,
    new_n17357_, new_n17358_, new_n17359_, new_n17360_, new_n17362_,
    new_n17363_, new_n17364_, new_n17365_, new_n17366_, new_n17367_,
    new_n17368_, new_n17369_, new_n17370_, new_n17371_, new_n17372_,
    new_n17373_, new_n17374_, new_n17375_, new_n17376_, new_n17377_,
    new_n17378_, new_n17380_, new_n17381_, new_n17382_, new_n17383_,
    new_n17384_, new_n17385_, new_n17386_, new_n17387_, new_n17388_,
    new_n17389_, new_n17390_, new_n17391_, new_n17392_, new_n17393_,
    new_n17394_, new_n17395_, new_n17396_, new_n17398_, new_n17399_,
    new_n17400_, new_n17401_, new_n17402_, new_n17403_, new_n17404_,
    new_n17405_, new_n17406_, new_n17407_, new_n17408_, new_n17409_,
    new_n17410_, new_n17411_, new_n17412_, new_n17413_, new_n17414_,
    new_n17415_, new_n17416_, new_n17417_, new_n17418_, new_n17420_,
    new_n17421_, new_n17422_, new_n17424_, new_n17425_, new_n17426_,
    new_n17428_, new_n17429_, new_n17430_, new_n17431_, new_n17432_,
    new_n17433_, new_n17434_, new_n17435_, new_n17436_, new_n17437_,
    new_n17438_, new_n17439_, new_n17440_, new_n17441_, new_n17442_,
    new_n17443_, new_n17444_, new_n17447_, new_n17448_, new_n17449_,
    new_n17451_, new_n17452_, new_n17453_, new_n17454_, new_n17455_,
    new_n17456_, new_n17457_, new_n17458_, new_n17459_, new_n17460_,
    new_n17461_, new_n17462_, new_n17463_, new_n17464_, new_n17465_,
    new_n17466_, new_n17467_, new_n17468_, new_n17469_, new_n17470_,
    new_n17471_, new_n17473_, new_n17474_, new_n17475_, new_n17477_,
    new_n17478_, new_n17479_, new_n17481_, new_n17482_, new_n17483_,
    new_n17485_, new_n17486_, new_n17487_, new_n17488_, new_n17489_,
    new_n17490_, new_n17491_, new_n17492_, new_n17493_, new_n17494_,
    new_n17495_, new_n17496_, new_n17497_, new_n17498_, new_n17499_,
    new_n17500_, new_n17501_, new_n17502_, new_n17503_, new_n17504_,
    new_n17505_, new_n17507_, new_n17508_, new_n17509_, new_n17511_,
    new_n17512_, new_n17513_, new_n17515_, new_n17516_, new_n17517_,
    new_n17518_, new_n17519_, new_n17520_, new_n17521_, new_n17522_,
    new_n17523_, new_n17524_, new_n17525_, new_n17526_, new_n17527_,
    new_n17528_, new_n17529_, new_n17530_, new_n17531_, new_n17532_,
    new_n17533_, new_n17534_, new_n17535_, new_n17537_, new_n17538_,
    new_n17539_, new_n17541_, new_n17542_, new_n17543_, new_n17545_,
    new_n17546_, new_n17547_, new_n17549_, new_n17550_, new_n17551_,
    new_n17553_, new_n17554_, new_n17555_, new_n17557_, new_n17558_,
    new_n17559_, new_n17561_, new_n17562_, new_n17563_, new_n17565_,
    new_n17566_, new_n17567_, new_n17569_, new_n17570_, new_n17571_,
    new_n17573_, new_n17574_, new_n17575_, new_n17577_, new_n17578_,
    new_n17579_, new_n17581_, new_n17582_, new_n17583_, new_n17585_,
    new_n17586_, new_n17587_, new_n17589_, new_n17590_, new_n17591_,
    new_n17593_, new_n17594_, new_n17595_, new_n17596_, new_n17597_,
    new_n17598_, new_n17599_, new_n17600_, new_n17601_, new_n17602_,
    new_n17603_, new_n17604_, new_n17605_, new_n17606_, new_n17607_,
    new_n17608_, new_n17609_, new_n17610_, new_n17611_, new_n17613_,
    new_n17614_, new_n17615_, new_n17616_, new_n17617_, new_n17618_,
    new_n17619_, new_n17620_, new_n17621_, new_n17622_, new_n17623_,
    new_n17624_, new_n17625_, new_n17626_, new_n17627_, new_n17628_,
    new_n17629_, new_n17630_, new_n17631_, new_n17633_, new_n17634_,
    new_n17635_, new_n17637_, new_n17638_, new_n17639_, new_n17641_,
    new_n17642_, new_n17643_, new_n17644_, new_n17645_, new_n17646_,
    new_n17647_, new_n17648_, new_n17649_, new_n17650_, new_n17651_,
    new_n17652_, new_n17653_, new_n17654_, new_n17655_, new_n17656_,
    new_n17657_, new_n17658_, new_n17659_, new_n17661_, new_n17662_,
    new_n17663_, new_n17664_, new_n17665_, new_n17666_, new_n17667_,
    new_n17668_, new_n17669_, new_n17670_, new_n17671_, new_n17672_,
    new_n17673_, new_n17674_, new_n17675_, new_n17676_, new_n17677_,
    new_n17678_, new_n17679_, new_n17681_, new_n17682_, new_n17683_,
    new_n17684_, new_n17685_, new_n17686_, new_n17687_, new_n17688_,
    new_n17689_, new_n17690_, new_n17691_, new_n17692_, new_n17693_,
    new_n17694_, new_n17695_, new_n17696_, new_n17697_, new_n17698_,
    new_n17699_, new_n17701_, new_n17702_, new_n17703_, new_n17704_,
    new_n17705_, new_n17706_, new_n17707_, new_n17708_, new_n17709_,
    new_n17710_, new_n17711_, new_n17712_, new_n17713_, new_n17714_,
    new_n17715_, new_n17716_, new_n17717_, new_n17718_, new_n17719_,
    new_n17720_, new_n17721_, new_n17723_, new_n17724_, new_n17725_,
    new_n17727_, new_n17728_, new_n17729_, new_n17730_, new_n17731_,
    new_n17732_, new_n17733_, new_n17734_, new_n17735_, new_n17736_,
    new_n17737_, new_n17738_, new_n17739_, new_n17740_, new_n17741_,
    new_n17742_, new_n17743_, new_n17744_, new_n17745_, new_n17747_,
    new_n17748_, new_n17749_, new_n17750_, new_n17751_, new_n17752_,
    new_n17753_, new_n17754_, new_n17755_, new_n17756_, new_n17757_,
    new_n17758_, new_n17759_, new_n17760_, new_n17761_, new_n17762_,
    new_n17763_, new_n17764_, new_n17765_, new_n17766_, new_n17767_,
    new_n17769_, new_n17770_, new_n17771_, new_n17772_, new_n17773_,
    new_n17774_, new_n17775_, new_n17776_, new_n17777_, new_n17778_,
    new_n17779_, new_n17780_, new_n17781_, new_n17782_, new_n17783_,
    new_n17784_, new_n17785_, new_n17786_, new_n17787_, new_n17789_,
    new_n17790_, new_n17791_, new_n17792_, new_n17793_, new_n17794_,
    new_n17795_, new_n17796_, new_n17797_, new_n17798_, new_n17799_,
    new_n17800_, new_n17801_, new_n17802_, new_n17803_, new_n17804_,
    new_n17805_, new_n17806_, new_n17807_, new_n17808_, new_n17809_,
    new_n17811_, new_n17812_, new_n17813_, new_n17814_, new_n17815_,
    new_n17816_, new_n17817_, new_n17818_, new_n17819_, new_n17820_,
    new_n17821_, new_n17822_, new_n17823_, new_n17824_, new_n17825_,
    new_n17826_, new_n17827_, new_n17828_, new_n17829_, new_n17830_,
    new_n17831_, new_n17833_, new_n17834_, new_n17835_, new_n17836_,
    new_n17837_, new_n17838_, new_n17839_, new_n17840_, new_n17841_,
    new_n17842_, new_n17843_, new_n17844_, new_n17845_, new_n17846_,
    new_n17847_, new_n17848_, new_n17849_, new_n17850_, new_n17851_,
    new_n17852_, new_n17853_, new_n17854_, new_n17855_, new_n17856_,
    new_n17857_, new_n17858_, new_n17859_, new_n17860_, new_n17861_,
    new_n17862_, new_n17863_, new_n17864_, new_n17865_, new_n17866_,
    new_n17867_, new_n17868_, new_n17869_, new_n17870_, new_n17871_,
    new_n17872_, new_n17873_, new_n17874_, new_n17875_, new_n17876_,
    new_n17877_, new_n17878_, new_n17879_, new_n17880_, new_n17882_,
    new_n17885_, new_n17886_, new_n17887_, new_n17888_, new_n17889_,
    new_n17890_, new_n17891_, new_n17892_, new_n17893_, new_n17894_,
    new_n17895_, new_n17896_, new_n17897_, new_n17898_, new_n17899_,
    new_n17900_, new_n17901_, new_n17902_, new_n17903_, new_n17904_,
    new_n17905_, new_n17907_, new_n17908_, new_n17909_, new_n17911_,
    new_n17912_, new_n17913_, new_n17915_, new_n17916_, new_n17917_,
    new_n17919_, new_n17920_, new_n17921_, new_n17923_, new_n17924_,
    new_n17925_, new_n17927_, new_n17928_, new_n17929_, new_n17931_,
    new_n17932_, new_n17933_, new_n17935_, new_n17936_, new_n17937_,
    new_n17939_, new_n17940_, new_n17941_, new_n17942_, new_n17943_,
    new_n17944_, new_n17945_, new_n17947_, new_n17948_, new_n17949_,
    new_n17951_, new_n17952_, new_n17953_, new_n17954_, new_n17955_,
    new_n17956_, new_n17957_, new_n17958_, new_n17959_, new_n17960_,
    new_n17961_, new_n17962_, new_n17963_, new_n17964_, new_n17965_,
    new_n17966_, new_n17967_, new_n17968_, new_n17969_, new_n17971_,
    new_n17972_, new_n17973_, new_n17975_, new_n17976_, new_n17977_,
    new_n17979_, new_n17980_, new_n17981_, new_n17983_, new_n17984_,
    new_n17985_, new_n17987_, new_n17988_, new_n17989_, new_n17992_,
    new_n17993_, new_n17994_, new_n17996_, new_n17997_, new_n17998_,
    new_n18000_, new_n18001_, new_n18002_, new_n18004_, new_n18005_,
    new_n18006_, new_n18008_, new_n18009_, new_n18010_, new_n18012_,
    new_n18013_, new_n18014_, new_n18016_, new_n18017_, new_n18018_,
    new_n18020_, new_n18021_, new_n18022_, new_n18023_, new_n18024_,
    new_n18026_, new_n18027_, new_n18028_, new_n18030_, new_n18031_,
    new_n18032_, new_n18034_, new_n18035_, new_n18036_, new_n18038_,
    new_n18039_, new_n18040_, new_n18042_, new_n18043_, new_n18044_,
    new_n18046_, new_n18047_, new_n18048_, new_n18050_, new_n18051_,
    new_n18052_, new_n18054_, new_n18055_, new_n18056_, new_n18058_,
    new_n18059_, new_n18060_, new_n18062_, new_n18063_, new_n18064_,
    new_n18066_, new_n18067_, new_n18068_, new_n18070_, new_n18071_,
    new_n18072_, new_n18074_, new_n18075_, new_n18076_, new_n18078_,
    new_n18079_, new_n18080_, new_n18082_, new_n18083_, new_n18084_,
    new_n18086_, new_n18087_, new_n18088_, new_n18090_, new_n18091_,
    new_n18092_, new_n18094_, new_n18095_, new_n18096_, new_n18098_,
    new_n18099_, new_n18100_, new_n18102_, new_n18103_, new_n18104_,
    new_n18106_, new_n18107_, new_n18108_, new_n18110_, new_n18111_,
    new_n18112_, new_n18113_, new_n18114_, new_n18115_, new_n18116_,
    new_n18117_, new_n18118_, new_n18120_, new_n18121_, new_n18122_,
    new_n18124_, new_n18125_, new_n18126_, new_n18127_, new_n18128_,
    new_n18129_, new_n18131_, new_n18132_, new_n18133_, new_n18135_,
    new_n18136_, new_n18137_, new_n18138_, new_n18139_, new_n18141_,
    new_n18142_, new_n18143_, new_n18145_, new_n18146_, new_n18147_,
    new_n18148_, new_n18149_, new_n18150_, new_n18151_, new_n18152_,
    new_n18153_, new_n18155_, new_n18156_, new_n18157_, new_n18159_,
    new_n18160_, new_n18161_, new_n18163_, new_n18164_, new_n18165_,
    new_n18166_, new_n18167_, new_n18168_, new_n18169_, new_n18173_,
    new_n18174_, new_n18176_, new_n18177_, new_n18179_, new_n18180_,
    new_n18182_, new_n18183_, new_n18185_, new_n18186_, new_n18188_,
    new_n18189_, new_n18191_, new_n18192_, new_n18194_, new_n18195_,
    new_n18197_, new_n18198_, new_n18200_, new_n18201_, new_n18203_,
    new_n18204_, new_n18206_, new_n18207_, new_n18209_, new_n18210_,
    new_n18211_, new_n18212_, new_n18214_, new_n18215_, new_n18217_,
    new_n18218_, new_n18219_, new_n18220_, new_n18221_, new_n18222_,
    new_n18223_, new_n18224_, new_n18225_, new_n18226_, new_n18228_,
    new_n18229_, new_n18231_, new_n18232_, new_n18234_, new_n18235_,
    new_n18237_, new_n18238_, new_n18240_, new_n18241_, new_n18242_,
    new_n18243_, new_n18244_, new_n18245_, new_n18247_, new_n18248_,
    new_n18250_, new_n18251_, new_n18253_, new_n18254_, new_n18256_,
    new_n18257_, new_n18259_, new_n18260_, new_n18262_, new_n18263_,
    new_n18265_, new_n18266_, new_n18268_, new_n18269_, new_n18271_,
    new_n18272_, new_n18274_, new_n18275_, new_n18277_, new_n18278_,
    new_n18280_, new_n18281_, new_n18283_, new_n18284_, new_n18286_,
    new_n18287_, new_n18289_, new_n18290_, new_n18291_, new_n18292_,
    new_n18293_, new_n18294_, new_n18296_, new_n18297_, new_n18298_,
    new_n18301_, new_n18302_, new_n18303_, new_n18305_, new_n18306_,
    new_n18307_, new_n18308_, new_n18309_, new_n18310_, new_n18311_,
    new_n18312_, new_n18313_, new_n18314_, new_n18315_, new_n18316_,
    new_n18317_, new_n18318_, new_n18319_, new_n18320_, new_n18321_,
    new_n18322_, new_n18323_, new_n18324_, new_n18325_, new_n18326_,
    new_n18327_, new_n18328_, new_n18330_, new_n18331_, new_n18332_,
    new_n18333_, new_n18334_, new_n18335_, new_n18336_, new_n18337_,
    new_n18338_, new_n18339_, new_n18340_, new_n18341_, new_n18342_,
    new_n18343_, new_n18344_, new_n18345_, new_n18346_, new_n18347_,
    new_n18348_, new_n18349_, new_n18350_, new_n18351_, new_n18352_,
    new_n18354_, new_n18355_, new_n18356_, new_n18357_, new_n18358_,
    new_n18359_, new_n18360_, new_n18361_, new_n18362_, new_n18363_,
    new_n18364_, new_n18365_, new_n18366_, new_n18367_, new_n18368_,
    new_n18369_, new_n18370_, new_n18371_, new_n18372_, new_n18373_,
    new_n18374_, new_n18375_, new_n18376_, new_n18378_, new_n18379_,
    new_n18380_, new_n18381_, new_n18382_, new_n18383_, new_n18384_,
    new_n18385_, new_n18386_, new_n18387_, new_n18388_, new_n18389_,
    new_n18390_, new_n18391_, new_n18392_, new_n18393_, new_n18394_,
    new_n18395_, new_n18396_, new_n18397_, new_n18398_, new_n18399_,
    new_n18400_, new_n18402_, new_n18403_, new_n18405_, new_n18406_,
    new_n18407_, new_n18409_, new_n18410_, new_n18412_, new_n18415_,
    new_n18416_, new_n18418_, new_n18419_, new_n18421_, new_n18422_,
    new_n18424_, new_n18425_, new_n18427_, new_n18428_, new_n18430_,
    new_n18431_, new_n18433_, new_n18434_, new_n18436_, new_n18437_,
    new_n18439_, new_n18440_, new_n18442_, new_n18443_, new_n18445_,
    new_n18446_, new_n18448_, new_n18449_, new_n18451_, new_n18452_,
    new_n18454_, new_n18455_, new_n18457_, new_n18458_, new_n18460_,
    new_n18461_, new_n18463_, new_n18464_, new_n18466_, new_n18467_,
    new_n18469_, new_n18470_, new_n18472_, new_n18473_, new_n18475_,
    new_n18476_, new_n18478_, new_n18479_, new_n18481_, new_n18482_,
    new_n18484_, new_n18485_, new_n18487_, new_n18488_, new_n18490_,
    new_n18491_, new_n18493_, new_n18494_, new_n18496_, new_n18497_,
    new_n18499_, new_n18500_, new_n18502_, new_n18503_, new_n18505_,
    new_n18506_, new_n18508_, new_n18509_, new_n18511_, new_n18512_,
    new_n18514_, new_n18515_, new_n18517_, new_n18518_, new_n18520_,
    new_n18521_, new_n18523_, new_n18524_, new_n18526_, new_n18527_,
    new_n18529_, new_n18530_, new_n18532_, new_n18533_, new_n18535_,
    new_n18536_, new_n18538_, new_n18539_, new_n18541_, new_n18542_,
    new_n18544_, new_n18545_, new_n18547_, new_n18548_, new_n18550_,
    new_n18551_, new_n18553_, new_n18554_, new_n18556_, new_n18557_,
    new_n18559_, new_n18560_, new_n18562_, new_n18563_, new_n18565_,
    new_n18566_, new_n18568_, new_n18569_, new_n18571_, new_n18572_,
    new_n18574_, new_n18575_, new_n18577_, new_n18578_, new_n18580_,
    new_n18581_, new_n18583_, new_n18584_, new_n18586_, new_n18587_,
    new_n18589_, new_n18590_, new_n18592_, new_n18593_, new_n18595_,
    new_n18596_, new_n18598_, new_n18599_, new_n18601_, new_n18602_,
    new_n18604_, new_n18605_, new_n18607_, new_n18608_, new_n18610_,
    new_n18611_, new_n18613_, new_n18614_, new_n18615_, new_n18616_,
    new_n18617_, new_n18618_, new_n18619_, new_n18620_, new_n18621_,
    new_n18623_, new_n18624_, new_n18626_, new_n18627_, new_n18629_,
    new_n18630_, new_n18632_, new_n18633_, new_n18635_, new_n18636_,
    new_n18638_, new_n18639_, new_n18641_, new_n18642_, new_n18644_,
    new_n18645_, new_n18647_, new_n18648_, new_n18650_, new_n18651_,
    new_n18653_, new_n18654_, new_n18656_, new_n18657_, new_n18659_,
    new_n18660_, new_n18662_, new_n18663_, new_n18665_, new_n18666_,
    new_n18668_, new_n18669_, new_n18671_, new_n18673_, new_n18674_,
    new_n18676_, new_n18677_, new_n18679_, new_n18680_, new_n18682_,
    new_n18683_, new_n18685_, new_n18686_, new_n18688_, new_n18689_,
    new_n18691_, new_n18692_, new_n18694_, new_n18695_, new_n18697_,
    new_n18698_, new_n18700_, new_n18701_, new_n18703_, new_n18704_,
    new_n18706_, new_n18707_, new_n18709_, new_n18710_, new_n18712_,
    new_n18713_, new_n18715_, new_n18716_, new_n18718_, new_n18719_,
    new_n18721_, new_n18722_, new_n18724_, new_n18725_, new_n18727_,
    new_n18728_, new_n18730_, new_n18731_, new_n18734_, new_n18735_,
    new_n18737_, new_n18738_, new_n18740_, new_n18741_, new_n18743_,
    new_n18745_, new_n18746_, li0000, li0001, li0002, li0003, li0004,
    li0005, li0006, li0007, li0008, li0009, li0010, li0011, li0012, li0013,
    li0014, li0015, li0016, li0017, li0018, li0019, li0020, li0021, li0022,
    li0023, li0024, li0025, li0026, li0027, li0028, li0029, li0030, li0031,
    li0032, li0033, li0034, li0035, li0036, li0037, li0038, li0039, li0040,
    li0041, li0042, li0043, li0044, li0045, li0046, li0047, li0048, li0049,
    li0050, li0051, li0052, li0053, li0054, li0055, li0056, li0057, li0058,
    li0059, li0060, li0061, li0062, li0063, li0064, li0065, li0066, li0067,
    li0068, li0069, li0070, li0071, li0072, li0073, li0074, li0075, li0076,
    li0077, li0078, li0079, li0080, li0081, li0082, li0083, li0084, li0085,
    li0086, li0087, li0088, li0089, li0090, li0091, li0092, li0093, li0094,
    li0095, li0096, li0097, li0098, li0099, li0100, li0101, li0102, li0103,
    li0104, li0105, li0106, li0107, li0108, li0109, li0110, li0111, li0112,
    li0113, li0114, li0115, li0116, li0117, li0118, li0119, li0120, li0121,
    li0122, li0123, li0124, li0125, li0126, li0127, li0128, li0129, li0130,
    li0131, li0132, li0133, li0134, li0135, li0136, li0137, li0138, li0139,
    li0140, li0141, li0142, li0143, li0144, li0145, li0146, li0147, li0148,
    li0149, li0150, li0151, li0152, li0153, li0154, li0155, li0156, li0157,
    li0158, li0159, li0160, li0161, li0162, li0163, li0164, li0165, li0166,
    li0167, li0168, li0169, li0170, li0171, li0172, li0173, li0174, li0175,
    li0176, li0177, li0178, li0179, li0180, li0181, li0182, li0183, li0184,
    li0185, li0186, li0187, li0188, li0189, li0190, li0191, li0192, li0193,
    li0194, li0195, li0196, li0197, li0198, li0199, li0200, li0201, li0202,
    li0203, li0204, li0205, li0206, li0207, li0208, li0209, li0210, li0211,
    li0212, li0213, li0214, li0215, li0216, li0217, li0218, li0219, li0220,
    li0221, li0222, li0223, li0224, li0225, li0226, li0227, li0228, li0229,
    li0230, li0231, li0232, li0233, li0234, li0235, li0236, li0237, li0238,
    li0239, li0240, li0241, li0242, li0243, li0244, li0245, li0246, li0247,
    li0248, li0249, li0250, li0251, li0252, li0253, li0254, li0255, li0256,
    li0257, li0258, li0259, li0260, li0261, li0262, li0263, li0264, li0265,
    li0266, li0267, li0268, li0269, li0270, li0271, li0272, li0273, li0274,
    li0275, li0276, li0277, li0278, li0279, li0280, li0281, li0282, li0283,
    li0284, li0285, li0286, li0287, li0288, li0289, li0290, li0291, li0292,
    li0293, li0294, li0295, li0296, li0297, li0298, li0299, li0300, li0301,
    li0302, li0303, li0304, li0305, li0306, li0307, li0308, li0309, li0310,
    li0311, li0312, li0313, li0314, li0315, li0316, li0317, li0318, li0319,
    li0320, li0321, li0322, li0323, li0324, li0325, li0326, li0327, li0328,
    li0329, li0330, li0331, li0332, li0333, li0334, li0335, li0336, li0337,
    li0338, li0339, li0340, li0341, li0342, li0343, li0344, li0345, li0346,
    li0347, li0348, li0349, li0350, li0351, li0352, li0353, li0354, li0355,
    li0356, li0357, li0358, li0359, li0360, li0361, li0362, li0363, li0364,
    li0365, li0366, li0367, li0368, li0369, li0370, li0371, li0372, li0373,
    li0374, li0375, li0376, li0377, li0378, li0379, li0380, li0381, li0382,
    li0383, li0384, li0385, li0386, li0387, li0388, li0389, li0390, li0391,
    li0392, li0393, li0394, li0395, li0396, li0397, li0398, li0399, li0400,
    li0401, li0402, li0403, li0404, li0405, li0406, li0407, li0408, li0409,
    li0410, li0411, li0412, li0413, li0414, li0415, li0416, li0417, li0418,
    li0419, li0420, li0421, li0422, li0423, li0424, li0425, li0426, li0427,
    li0428, li0429, li0430, li0431, li0432, li0433, li0434, li0435, li0436,
    li0437, li0438, li0439, li0440, li0441, li0442, li0443, li0444, li0445,
    li0446, li0447, li0448, li0449, li0450, li0451, li0452, li0453, li0454,
    li0455, li0456, li0457, li0458, li0459, li0460, li0461, li0462, li0463,
    li0464, li0465, li0466, li0467, li0468, li0469, li0470, li0471, li0472,
    li0473, li0474, li0475, li0476, li0477, li0478, li0479, li0480, li0481,
    li0482, li0483, li0484, li0485, li0486, li0487, li0488, li0489, li0490,
    li0491, li0492, li0493, li0494, li0495, li0496, li0497, li0498, li0499,
    li0500, li0501, li0502, li0503, li0504, li0505, li0506, li0507, li0508,
    li0509, li0510, li0511, li0512, li0513, li0514, li0515, li0516, li0517,
    li0518, li0519, li0520, li0521, li0522, li0523, li0524, li0525, li0526,
    li0527, li0528, li0529, li0530, li0531, li0532, li0533, li0534, li0535,
    li0536, li0537, li0538, li0539, li0540, li0541, li0542, li0543, li0544,
    li0545, li0546, li0547, li0548, li0549, li0550, li0551, li0552, li0553,
    li0554, li0555, li0556, li0557, li0558, li0559, li0560, li0561, li0562,
    li0563, li0564, li0565, li0566, li0567, li0568, li0569, li0570, li0571,
    li0572, li0573, li0574, li0575, li0576, li0577, li0578, li0579, li0580,
    li0581, li0582, li0583, li0584, li0585, li0586, li0587, li0588, li0589,
    li0590, li0591, li0592, li0593, li0594, li0595, li0596, li0597, li0598,
    li0599, li0600, li0601, li0602, li0603, li0604, li0605, li0606, li0607,
    li0608, li0609, li0610, li0611, li0612, li0613, li0614, li0615, li0616,
    li0617, li0618, li0619, li0620, li0621, li0622, li0623, li0624, li0625,
    li0626, li0627, li0628, li0629, li0630, li0631, li0632, li0633, li0634,
    li0635, li0636, li0637, li0638, li0639, li0640, li0641, li0642, li0643,
    li0644, li0645, li0646, li0647, li0648, li0649, li0650, li0651, li0652,
    li0653, li0654, li0655, li0656, li0657, li0658, li0659, li0660, li0661,
    li0662, li0663, li0664, li0665, li0666, li0667, li0668, li0669, li0670,
    li0671, li0672, li0673, li0674, li0675, li0676, li0677, li0678, li0679,
    li0680, li0681, li0682, li0683, li0684, li0685, li0686, li0687, li0688,
    li0689, li0690, li0691, li0692, li0693, li0694, li0695, li0696, li0697,
    li0698, li0699, li0700, li0701, li0702, li0703, li0704, li0705, li0706,
    li0707, li0708, li0709, li0710, li0711, li0712, li0713, li0714, li0715,
    li0716, li0717, li0718, li0719, li0720, li0721, li0722, li0723, li0724,
    li0725, li0726, li0727, li0728, li0729, li0730, li0731, li0732, li0733,
    li0734, li0735, li0736, li0737, li0738, li0739, li0740, li0741, li0742,
    li0743, li0744, li0745, li0746, li0747, li0748, li0749, li0750, li0751,
    li0752, li0753, li0754, li0755, li0756, li0757, li0758, li0759, li0760,
    li0761, li0762, li0763, li0764, li0765, li0766, li0767, li0768, li0769,
    li0770, li0771, li0772, li0773, li0774, li0775, li0776, li0777, li0778,
    li0779, li0780, li0781, li0782, li0783, li0784, li0785, li0786, li0787,
    li0788, li0789, li0790, li0791, li0792, li0793, li0794, li0795, li0796,
    li0797, li0798, li0799, li0800, li0801, li0802, li0803, li0804, li0805,
    li0806, li0807, li0808, li0809, li0810, li0811, li0812, li0813, li0814,
    li0815, li0816, li0817, li0818, li0819, li0820, li0821, li0822, li0823,
    li0824, li0825, li0826, li0827, li0828, li0829, li0830, li0831, li0832,
    li0833, li0834, li0835, li0836, li0837, li0838, li0839, li0840, li0841,
    li0842, li0843, li0844, li0845, li0846, li0847, li0848, li0849, li0850,
    li0851, li0852, li0853, li0854, li0855, li0856, li0857, li0858, li0859,
    li0860, li0861, li0862, li0863, li0864, li0865, li0866, li0867, li0868,
    li0869, li0870, li0871, li0872, li0873, li0874, li0875, li0876, li0877,
    li0878, li0879, li0880, li0881, li0882, li0883, li0884, li0885, li0886,
    li0887, li0888, li0889, li0890, li0891, li0892, li0893, li0894, li0895,
    li0896, li0897, li0898, li0899, li0900, li0901, li0902, li0903, li0904,
    li0905, li0906, li0907, li0908, li0909, li0910, li0911, li0912, li0913,
    li0914, li0915, li0916, li0917, li0918, li0919, li0920, li0921, li0922,
    li0923, li0924, li0925, li0926, li0927, li0928, li0929, li0930, li0931,
    li0932, li0933, li0934, li0935, li0936, li0937, li0938, li0939, li0940,
    li0941, li0942, li0943, li0944, li0945, li0946, li0947, li0948, li0949,
    li0950, li0951, li0952, li0953, li0954, li0955, li0956, li0957, li0958,
    li0959, li0960, li0961, li0962, li0963, li0964, li0965, li0966, li0967,
    li0968, li0969, li0970, li0971, li0972, li0973, li0974, li0975, li0976,
    li0977, li0978, li0979, li0980, li0981, li0982, li0983, li0984, li0985,
    li0986, li0987, li0988, li0989, li0990, li0991, li0992, li0993, li0994,
    li0995, li0996, li0997, li0998, li0999, li1000, li1001, li1002, li1003,
    li1004, li1005, li1006, li1007, li1008, li1009, li1010, li1011, li1012,
    li1013, li1014, li1015, li1016, li1017, li1018, li1019, li1020, li1021,
    li1022, li1023, li1024, li1025, li1026, li1027, li1028, li1029, li1030,
    li1031, li1032, li1033, li1034, li1035, li1036, li1037, li1038, li1039,
    li1040, li1041, li1042, li1043, li1044, li1045, li1046, li1047, li1048,
    li1049, li1050, li1051, li1052, li1053, li1054, li1055, li1056, li1057,
    li1058, li1059, li1060, li1061, li1062, li1063, li1064, li1065, li1066,
    li1067, li1068, li1069, li1070, li1071, li1072, li1073, li1074, li1075,
    li1076, li1077, li1078, li1079, li1080, li1081, li1082;
  assign new_n3518_ = ~lo0057 & ~lo0059;
  assign new_n3519_ = ~lo0055 & ~lo0299;
  assign new_n3520_ = ~lo0056 & ~lo0062;
  assign new_n3521_ = new_n3518_ & new_n3519_;
  assign new_n3522_ = new_n3520_ & new_n3521_;
  assign new_n3523_ = lo0153 & ~new_n3522_;
  assign new_n3524_ = lo0175 & new_n3522_;
  assign new_n3525_ = ~new_n3523_ & ~new_n3524_;
  assign new_n3526_ = ~lo0035 & ~lo0070;
  assign new_n3527_ = ~lo0049 & ~lo0076;
  assign new_n3528_ = ~lo0075 & ~lo0094;
  assign new_n3529_ = new_n3526_ & new_n3527_;
  assign new_n3530_ = new_n3528_ & new_n3529_;
  assign new_n3531_ = lo0089 & new_n3530_;
  assign new_n3532_ = ~lo0095 & ~lo0097;
  assign new_n3533_ = ~lo0074 & ~lo0096;
  assign new_n3534_ = new_n3532_ & new_n3533_;
  assign new_n3535_ = ~lo0032 & ~lo0038;
  assign new_n3536_ = ~lo0050 & ~lo0100;
  assign new_n3537_ = new_n3535_ & new_n3536_;
  assign new_n3538_ = new_n3534_ & new_n3537_;
  assign new_n3539_ = ~lo0108 & new_n3538_;
  assign new_n3540_ = ~lo0039 & ~lo0048;
  assign new_n3541_ = ~lo0087 & ~lo0111;
  assign new_n3542_ = ~lo0072 & ~lo0103;
  assign new_n3543_ = new_n3541_ & new_n3542_;
  assign new_n3544_ = ~lo0088 & ~lo0104;
  assign new_n3545_ = ~lo0047 & ~lo0110;
  assign new_n3546_ = new_n3544_ & new_n3545_;
  assign new_n3547_ = new_n3543_ & new_n3546_;
  assign new_n3548_ = ~lo0073 & ~lo0090;
  assign new_n3549_ = ~lo0036 & ~lo0091;
  assign new_n3550_ = new_n3548_ & new_n3549_;
  assign new_n3551_ = ~lo0092 & ~lo0093;
  assign new_n3552_ = ~lo0058 & ~lo0098;
  assign new_n3553_ = new_n3551_ & new_n3552_;
  assign new_n3554_ = new_n3550_ & new_n3553_;
  assign new_n3555_ = new_n3540_ & new_n3547_;
  assign new_n3556_ = new_n3554_ & new_n3555_;
  assign new_n3557_ = ~lo0066 & ~lo0082;
  assign new_n3558_ = ~lo0051 & ~lo0084;
  assign new_n3559_ = new_n3557_ & new_n3558_;
  assign new_n3560_ = ~lo0040 & ~lo0081;
  assign new_n3561_ = ~lo0068 & ~lo0102;
  assign new_n3562_ = new_n3560_ & new_n3561_;
  assign new_n3563_ = new_n3559_ & new_n3562_;
  assign new_n3564_ = ~lo0077 & ~lo0086;
  assign new_n3565_ = ~lo0069 & ~lo0109;
  assign new_n3566_ = new_n3564_ & new_n3565_;
  assign new_n3567_ = ~lo0067 & ~lo0071;
  assign new_n3568_ = ~lo0083 & ~lo0085;
  assign new_n3569_ = new_n3567_ & new_n3568_;
  assign new_n3570_ = new_n3563_ & new_n3566_;
  assign new_n3571_ = new_n3569_ & new_n3570_;
  assign new_n3572_ = ~lo0045 & ~lo0053;
  assign new_n3573_ = ~lo0054 & ~lo0106;
  assign new_n3574_ = new_n3572_ & new_n3573_;
  assign new_n3575_ = ~lo0055 & ~lo0057;
  assign new_n3576_ = new_n3520_ & new_n3575_;
  assign new_n3577_ = new_n3574_ & new_n3576_;
  assign new_n3578_ = ~lo0064 & ~lo0065;
  assign new_n3579_ = ~lo0063 & ~lo0107;
  assign new_n3580_ = new_n3578_ & new_n3579_;
  assign new_n3581_ = ~lo0046 & ~lo0061;
  assign new_n3582_ = ~lo0059 & ~lo0060;
  assign new_n3583_ = new_n3581_ & new_n3582_;
  assign new_n3584_ = new_n3580_ & new_n3583_;
  assign new_n3585_ = new_n3577_ & new_n3584_;
  assign new_n3586_ = new_n3556_ & new_n3571_;
  assign new_n3587_ = new_n3585_ & new_n3586_;
  assign new_n3588_ = new_n3539_ & new_n3587_;
  assign new_n3589_ = new_n3531_ & new_n3588_;
  assign new_n3590_ = new_n3527_ & new_n3528_;
  assign new_n3591_ = lo0070 & new_n3590_;
  assign new_n3592_ = ~lo0089 & ~lo0108;
  assign new_n3593_ = new_n3591_ & new_n3592_;
  assign new_n3594_ = ~lo0035 & new_n3593_;
  assign new_n3595_ = new_n3537_ & new_n3587_;
  assign new_n3596_ = new_n3534_ & new_n3595_;
  assign new_n3597_ = new_n3594_ & new_n3596_;
  assign new_n3598_ = ~new_n3589_ & ~new_n3597_;
  assign new_n3599_ = lo0287 & ~new_n3598_;
  assign new_n3600_ = ~lo0287 & lo0332;
  assign new_n3601_ = ~new_n3599_ & ~new_n3600_;
  assign new_n3602_ = new_n3547_ & new_n3554_;
  assign new_n3603_ = new_n3571_ & new_n3602_;
  assign new_n3604_ = new_n3526_ & new_n3592_;
  assign new_n3605_ = new_n3534_ & new_n3604_;
  assign new_n3606_ = new_n3536_ & new_n3590_;
  assign new_n3607_ = new_n3535_ & new_n3606_;
  assign new_n3608_ = new_n3605_ & new_n3607_;
  assign new_n3609_ = new_n3585_ & new_n3603_;
  assign new_n3610_ = new_n3608_ & new_n3609_;
  assign new_n3611_ = lo0039 & ~lo0048;
  assign new_n3612_ = new_n3610_ & new_n3611_;
  assign new_n3613_ = ~new_n3589_ & ~new_n3612_;
  assign new_n3614_ = ~new_n3601_ & ~new_n3613_;
  assign new_n3615_ = ~lo0032 & new_n3606_;
  assign new_n3616_ = lo0038 & new_n3605_;
  assign new_n3617_ = new_n3615_ & new_n3616_;
  assign new_n3618_ = new_n3587_ & new_n3617_;
  assign new_n3619_ = ~lo0061 & new_n3580_;
  assign new_n3620_ = lo0046 & new_n3582_;
  assign new_n3621_ = new_n3608_ & new_n3619_;
  assign new_n3622_ = new_n3620_ & new_n3621_;
  assign new_n3623_ = new_n3540_ & new_n3577_;
  assign new_n3624_ = new_n3622_ & new_n3623_;
  assign new_n3625_ = new_n3603_ & new_n3624_;
  assign new_n3626_ = ~new_n3618_ & ~new_n3625_;
  assign new_n3627_ = new_n3613_ & ~new_n3626_;
  assign new_n3628_ = new_n3598_ & new_n3627_;
  assign new_n3629_ = lo0332 & new_n3613_;
  assign new_n3630_ = ~new_n3598_ & new_n3629_;
  assign new_n3631_ = lo0152 & ~new_n3522_;
  assign new_n3632_ = lo0174 & new_n3522_;
  assign new_n3633_ = ~new_n3631_ & ~new_n3632_;
  assign new_n3634_ = ~lo0057 & new_n3520_;
  assign new_n3635_ = new_n3519_ & new_n3634_;
  assign new_n3636_ = ~lo0059 & new_n3635_;
  assign new_n3637_ = lo0144 & new_n3636_;
  assign new_n3638_ = lo0161 & ~new_n3522_;
  assign new_n3639_ = ~new_n3637_ & ~new_n3638_;
  assign new_n3640_ = new_n3633_ & new_n3639_;
  assign new_n3641_ = ~lo0332 & ~lo0468;
  assign new_n3642_ = lo0232 & new_n3641_;
  assign new_n3643_ = lo0189 & new_n3636_;
  assign new_n3644_ = lo0166 & ~new_n3636_;
  assign new_n3645_ = ~new_n3643_ & ~new_n3644_;
  assign new_n3646_ = new_n3642_ & new_n3645_;
  assign new_n3647_ = new_n3640_ & new_n3646_;
  assign new_n3648_ = ~new_n3614_ & ~new_n3628_;
  assign new_n3649_ = ~new_n3630_ & new_n3648_;
  assign new_n3650_ = new_n3647_ & new_n3649_;
  assign new_n3651_ = lo0142 & new_n3522_;
  assign new_n3652_ = lo0146 & ~new_n3522_;
  assign new_n3653_ = ~new_n3651_ & ~new_n3652_;
  assign new_n3654_ = new_n3640_ & new_n3645_;
  assign new_n3655_ = new_n3653_ & ~new_n3654_;
  assign new_n3656_ = ~lo0115 & ~lo0116;
  assign new_n3657_ = ~lo0099 & ~lo0113;
  assign new_n3658_ = new_n3656_ & new_n3657_;
  assign new_n3659_ = ~lo0044 & new_n3658_;
  assign new_n3660_ = ~lo0042 & ~lo0043;
  assign new_n3661_ = ~lo0041 & new_n3660_;
  assign new_n3662_ = ~lo0052 & new_n3661_;
  assign new_n3663_ = ~lo0114 & new_n3662_;
  assign new_n3664_ = ~lo0101 & new_n3663_;
  assign li0901 = ~new_n3659_ | ~new_n3664_;
  assign new_n3666_ = ~lo0683 & li0901;
  assign new_n3667_ = ~new_n3650_ & new_n3655_;
  assign new_n3668_ = new_n3666_ & new_n3667_;
  assign new_n3669_ = lo0252 & ~new_n3655_;
  assign new_n3670_ = ~lo0250 & new_n3655_;
  assign new_n3671_ = lo0129 & ~new_n3670_;
  assign new_n3672_ = pi002 & lo0957;
  assign new_n3673_ = pi003 & pi004;
  assign new_n3674_ = ~lo0833 & new_n3672_;
  assign li0950 = new_n3673_ & new_n3674_;
  assign li0982 = pi003 & lo0824;
  assign new_n3677_ = ~lo0950 & ~li0950;
  assign new_n3678_ = li0982 & new_n3677_;
  assign new_n3679_ = ~pi002 & pi004;
  assign new_n3680_ = pi003 & lo0829;
  assign li0951 = ~new_n3679_ & new_n3680_;
  assign new_n3682_ = ~lo0950 & li0951;
  assign li0683 = ~li0950 & new_n3682_;
  assign li0793 = ~new_n3678_ & ~li0683;
  assign new_n3685_ = pi003 & ~pi004;
  assign li0583 = ~li0793 & new_n3685_;
  assign new_n3687_ = new_n3670_ & ~li0583;
  assign new_n3688_ = ~lo0252 & ~new_n3655_;
  assign new_n3689_ = ~new_n3671_ & ~new_n3687_;
  assign new_n3690_ = ~new_n3688_ & ~new_n3689_;
  assign new_n3691_ = ~new_n3668_ & new_n3669_;
  assign new_n3692_ = new_n3690_ & ~new_n3691_;
  assign new_n3693_ = ~new_n3669_ & ~new_n3689_;
  assign new_n3694_ = new_n3688_ & new_n3693_;
  assign new_n3695_ = lo0100 & new_n3590_;
  assign new_n3696_ = ~lo0050 & new_n3695_;
  assign new_n3697_ = new_n3587_ & new_n3605_;
  assign new_n3698_ = new_n3535_ & new_n3697_;
  assign new_n3699_ = new_n3696_ & new_n3698_;
  assign new_n3700_ = ~new_n3692_ & ~new_n3694_;
  assign new_n3701_ = new_n3699_ & ~new_n3700_;
  assign new_n3702_ = lo0094 & new_n3527_;
  assign new_n3703_ = ~lo0075 & new_n3702_;
  assign new_n3704_ = new_n3537_ & new_n3697_;
  assign new_n3705_ = new_n3703_ & new_n3704_;
  assign new_n3706_ = new_n3689_ & new_n3699_;
  assign new_n3707_ = ~new_n3669_ & new_n3706_;
  assign new_n3708_ = new_n3577_ & new_n3583_;
  assign new_n3709_ = new_n3540_ & new_n3603_;
  assign new_n3710_ = new_n3708_ & new_n3709_;
  assign new_n3711_ = new_n3608_ & new_n3710_;
  assign new_n3712_ = lo0064 & ~lo0065;
  assign new_n3713_ = new_n3579_ & new_n3711_;
  assign new_n3714_ = new_n3712_ & new_n3713_;
  assign new_n3715_ = ~new_n3707_ & ~new_n3714_;
  assign new_n3716_ = new_n3562_ & new_n3566_;
  assign new_n3717_ = ~lo0066 & new_n3569_;
  assign new_n3718_ = new_n3716_ & new_n3717_;
  assign new_n3719_ = new_n3558_ & new_n3718_;
  assign new_n3720_ = lo0082 & new_n3719_;
  assign new_n3721_ = new_n3585_ & new_n3608_;
  assign new_n3722_ = new_n3556_ & new_n3721_;
  assign new_n3723_ = new_n3720_ & new_n3722_;
  assign new_n3724_ = ~lo0039 & lo0048;
  assign new_n3725_ = new_n3610_ & new_n3724_;
  assign new_n3726_ = ~new_n3723_ & ~new_n3725_;
  assign new_n3727_ = ~new_n3701_ & ~new_n3705_;
  assign new_n3728_ = new_n3715_ & new_n3727_;
  assign new_n3729_ = new_n3726_ & new_n3728_;
  assign new_n3730_ = new_n3577_ & new_n3709_;
  assign new_n3731_ = lo0061 & new_n3580_;
  assign new_n3732_ = ~lo0046 & new_n3582_;
  assign new_n3733_ = new_n3608_ & new_n3730_;
  assign new_n3734_ = new_n3731_ & new_n3733_;
  assign new_n3735_ = new_n3732_ & new_n3734_;
  assign new_n3736_ = ~lo0063 & lo0107;
  assign new_n3737_ = new_n3578_ & new_n3583_;
  assign new_n3738_ = new_n3733_ & new_n3736_;
  assign new_n3739_ = new_n3737_ & new_n3738_;
  assign new_n3740_ = ~new_n3735_ & ~new_n3739_;
  assign new_n3741_ = new_n3559_ & new_n3566_;
  assign new_n3742_ = new_n3561_ & new_n3569_;
  assign new_n3743_ = new_n3741_ & new_n3742_;
  assign new_n3744_ = ~lo0040 & new_n3743_;
  assign new_n3745_ = lo0081 & new_n3744_;
  assign new_n3746_ = new_n3722_ & new_n3745_;
  assign new_n3747_ = new_n3540_ & new_n3571_;
  assign new_n3748_ = new_n3721_ & new_n3747_;
  assign new_n3749_ = lo0036 & new_n3548_;
  assign new_n3750_ = ~lo0091 & new_n3553_;
  assign new_n3751_ = new_n3547_ & new_n3748_;
  assign new_n3752_ = new_n3749_ & new_n3751_;
  assign new_n3753_ = new_n3750_ & new_n3752_;
  assign new_n3754_ = new_n3740_ & ~new_n3746_;
  assign new_n3755_ = ~new_n3753_ & new_n3754_;
  assign new_n3756_ = new_n3613_ & new_n3755_;
  assign new_n3757_ = new_n3574_ & new_n3709_;
  assign new_n3758_ = new_n3583_ & new_n3757_;
  assign new_n3759_ = new_n3575_ & new_n3580_;
  assign new_n3760_ = ~lo0056 & lo0062;
  assign new_n3761_ = new_n3758_ & new_n3759_;
  assign new_n3762_ = new_n3608_ & new_n3761_;
  assign new_n3763_ = new_n3760_ & new_n3762_;
  assign new_n3764_ = new_n3546_ & new_n3550_;
  assign new_n3765_ = ~lo0111 & new_n3553_;
  assign new_n3766_ = lo0087 & new_n3542_;
  assign new_n3767_ = new_n3764_ & new_n3765_;
  assign new_n3768_ = new_n3766_ & new_n3767_;
  assign new_n3769_ = new_n3748_ & new_n3768_;
  assign new_n3770_ = ~new_n3763_ & ~new_n3769_;
  assign new_n3771_ = ~lo0081 & new_n3743_;
  assign new_n3772_ = lo0040 & new_n3722_;
  assign new_n3773_ = new_n3771_ & new_n3772_;
  assign new_n3774_ = new_n3770_ & ~new_n3773_;
  assign new_n3775_ = lo0076 & new_n3528_;
  assign new_n3776_ = ~lo0049 & new_n3775_;
  assign new_n3777_ = new_n3704_ & new_n3776_;
  assign new_n3778_ = lo0050 & ~lo0100;
  assign new_n3779_ = new_n3590_ & new_n3778_;
  assign new_n3780_ = new_n3698_ & new_n3779_;
  assign new_n3781_ = ~lo0059 & lo0060;
  assign new_n3782_ = new_n3709_ & new_n3781_;
  assign new_n3783_ = new_n3580_ & new_n3581_;
  assign new_n3784_ = new_n3608_ & new_n3782_;
  assign new_n3785_ = new_n3783_ & new_n3784_;
  assign new_n3786_ = new_n3577_ & new_n3785_;
  assign new_n3787_ = new_n3774_ & ~new_n3777_;
  assign new_n3788_ = ~new_n3780_ & new_n3787_;
  assign new_n3789_ = ~new_n3786_ & new_n3788_;
  assign new_n3790_ = new_n3564_ & new_n3569_;
  assign new_n3791_ = new_n3563_ & new_n3790_;
  assign new_n3792_ = ~lo0109 & new_n3791_;
  assign new_n3793_ = lo0069 & new_n3792_;
  assign new_n3794_ = new_n3722_ & new_n3793_;
  assign new_n3795_ = lo0086 & new_n3569_;
  assign new_n3796_ = new_n3563_ & new_n3795_;
  assign new_n3797_ = new_n3565_ & new_n3796_;
  assign new_n3798_ = ~lo0077 & new_n3797_;
  assign new_n3799_ = new_n3722_ & new_n3798_;
  assign new_n3800_ = ~new_n3794_ & ~new_n3799_;
  assign new_n3801_ = new_n3789_ & new_n3800_;
  assign new_n3802_ = ~lo0035 & new_n3591_;
  assign new_n3803_ = new_n3596_ & new_n3802_;
  assign new_n3804_ = new_n3592_ & new_n3803_;
  assign new_n3805_ = ~lo0074 & new_n3590_;
  assign new_n3806_ = lo0096 & new_n3805_;
  assign new_n3807_ = new_n3537_ & new_n3604_;
  assign new_n3808_ = new_n3587_ & new_n3807_;
  assign new_n3809_ = new_n3532_ & new_n3808_;
  assign new_n3810_ = new_n3806_ & new_n3809_;
  assign new_n3811_ = ~lo0072 & lo0103;
  assign new_n3812_ = new_n3764_ & new_n3811_;
  assign new_n3813_ = new_n3541_ & new_n3553_;
  assign new_n3814_ = new_n3748_ & new_n3812_;
  assign new_n3815_ = new_n3813_ & new_n3814_;
  assign new_n3816_ = lo0049 & new_n3534_;
  assign new_n3817_ = new_n3587_ & new_n3816_;
  assign new_n3818_ = new_n3528_ & new_n3817_;
  assign new_n3819_ = ~lo0076 & new_n3818_;
  assign new_n3820_ = new_n3807_ & new_n3819_;
  assign new_n3821_ = ~new_n3804_ & ~new_n3810_;
  assign new_n3822_ = ~new_n3815_ & new_n3821_;
  assign new_n3823_ = ~new_n3820_ & new_n3822_;
  assign new_n3824_ = lo0068 & new_n3569_;
  assign new_n3825_ = ~lo0102 & new_n3560_;
  assign new_n3826_ = new_n3722_ & new_n3824_;
  assign new_n3827_ = new_n3741_ & new_n3826_;
  assign new_n3828_ = new_n3825_ & new_n3827_;
  assign new_n3829_ = new_n3543_ & new_n3550_;
  assign new_n3830_ = new_n3545_ & new_n3553_;
  assign new_n3831_ = new_n3829_ & new_n3830_;
  assign new_n3832_ = ~lo0104 & new_n3831_;
  assign new_n3833_ = lo0088 & new_n3748_;
  assign new_n3834_ = new_n3832_ & new_n3833_;
  assign new_n3835_ = new_n3569_ & new_n3608_;
  assign new_n3836_ = new_n3556_ & new_n3585_;
  assign new_n3837_ = ~lo0051 & lo0084;
  assign new_n3838_ = new_n3557_ & new_n3837_;
  assign new_n3839_ = new_n3835_ & new_n3836_;
  assign new_n3840_ = new_n3716_ & new_n3839_;
  assign new_n3841_ = new_n3838_ & new_n3840_;
  assign new_n3842_ = ~lo0082 & new_n3558_;
  assign new_n3843_ = new_n3716_ & new_n3842_;
  assign new_n3844_ = lo0066 & new_n3843_;
  assign new_n3845_ = new_n3569_ & new_n3844_;
  assign new_n3846_ = new_n3722_ & new_n3845_;
  assign new_n3847_ = ~new_n3841_ & ~new_n3846_;
  assign new_n3848_ = ~new_n3828_ & ~new_n3834_;
  assign new_n3849_ = new_n3847_ & new_n3848_;
  assign new_n3850_ = new_n3823_ & new_n3849_;
  assign new_n3851_ = ~lo0073 & lo0090;
  assign new_n3852_ = new_n3608_ & new_n3851_;
  assign new_n3853_ = new_n3549_ & new_n3553_;
  assign new_n3854_ = new_n3547_ & new_n3853_;
  assign new_n3855_ = new_n3585_ & new_n3854_;
  assign new_n3856_ = new_n3747_ & new_n3852_;
  assign new_n3857_ = new_n3855_ & new_n3856_;
  assign new_n3858_ = new_n3550_ & new_n3552_;
  assign new_n3859_ = new_n3547_ & new_n3858_;
  assign new_n3860_ = lo0093 & new_n3859_;
  assign new_n3861_ = ~lo0092 & new_n3860_;
  assign new_n3862_ = new_n3748_ & new_n3861_;
  assign new_n3863_ = ~new_n3857_ & ~new_n3862_;
  assign new_n3864_ = ~lo0070 & new_n3590_;
  assign new_n3865_ = new_n3592_ & new_n3864_;
  assign new_n3866_ = lo0035 & new_n3865_;
  assign new_n3867_ = new_n3596_ & new_n3866_;
  assign new_n3868_ = lo0073 & ~lo0090;
  assign new_n3869_ = new_n3751_ & new_n3853_;
  assign new_n3870_ = new_n3868_ & new_n3869_;
  assign new_n3871_ = ~new_n3867_ & ~new_n3870_;
  assign new_n3872_ = new_n3863_ & new_n3871_;
  assign new_n3873_ = new_n3576_ & new_n3583_;
  assign new_n3874_ = new_n3709_ & new_n3873_;
  assign new_n3875_ = ~lo0053 & new_n3580_;
  assign new_n3876_ = lo0045 & new_n3573_;
  assign new_n3877_ = new_n3608_ & new_n3874_;
  assign new_n3878_ = new_n3875_ & new_n3877_;
  assign new_n3879_ = new_n3876_ & new_n3878_;
  assign new_n3880_ = new_n3872_ & ~new_n3879_;
  assign new_n3881_ = new_n3756_ & new_n3801_;
  assign new_n3882_ = new_n3850_ & new_n3881_;
  assign new_n3883_ = new_n3880_ & new_n3882_;
  assign new_n3884_ = lo0058 & new_n3550_;
  assign new_n3885_ = new_n3547_ & new_n3884_;
  assign new_n3886_ = ~lo0098 & new_n3885_;
  assign new_n3887_ = new_n3551_ & new_n3886_;
  assign new_n3888_ = new_n3748_ & new_n3887_;
  assign new_n3889_ = ~lo0088 & new_n3831_;
  assign new_n3890_ = lo0104 & new_n3889_;
  assign new_n3891_ = new_n3748_ & new_n3890_;
  assign new_n3892_ = ~new_n3888_ & ~new_n3891_;
  assign new_n3893_ = new_n3608_ & new_n3836_;
  assign new_n3894_ = new_n3566_ & new_n3893_;
  assign new_n3895_ = new_n3563_ & new_n3894_;
  assign new_n3896_ = ~lo0071 & new_n3895_;
  assign new_n3897_ = new_n3568_ & new_n3896_;
  assign new_n3898_ = lo0067 & new_n3897_;
  assign new_n3899_ = lo0083 & new_n3566_;
  assign new_n3900_ = new_n3563_ & new_n3567_;
  assign new_n3901_ = ~lo0085 & new_n3900_;
  assign new_n3902_ = new_n3722_ & new_n3899_;
  assign new_n3903_ = new_n3901_ & new_n3902_;
  assign new_n3904_ = ~new_n3898_ & ~new_n3903_;
  assign new_n3905_ = ~lo0067 & lo0071;
  assign new_n3906_ = new_n3568_ & new_n3905_;
  assign new_n3907_ = new_n3895_ & new_n3906_;
  assign new_n3908_ = new_n3556_ & new_n3608_;
  assign new_n3909_ = new_n3585_ & new_n3908_;
  assign new_n3910_ = lo0085 & new_n3567_;
  assign new_n3911_ = new_n3563_ & new_n3910_;
  assign new_n3912_ = ~lo0083 & new_n3566_;
  assign new_n3913_ = new_n3909_ & new_n3911_;
  assign new_n3914_ = new_n3912_ & new_n3913_;
  assign new_n3915_ = ~new_n3907_ & ~new_n3914_;
  assign new_n3916_ = new_n3904_ & new_n3915_;
  assign new_n3917_ = new_n3892_ & new_n3916_;
  assign new_n3918_ = new_n3608_ & new_n3708_;
  assign li0893 = lo0064 | ~new_n3579_;
  assign new_n3920_ = new_n3709_ & ~li0893;
  assign new_n3921_ = lo0065 & new_n3920_;
  assign new_n3922_ = new_n3918_ & new_n3921_;
  assign new_n3923_ = ~lo0228 & ~new_n3922_;
  assign new_n3924_ = new_n3917_ & new_n3923_;
  assign new_n3925_ = lo0063 & ~lo0107;
  assign new_n3926_ = new_n3733_ & new_n3737_;
  assign new_n3927_ = new_n3925_ & new_n3926_;
  assign new_n3928_ = lo0056 & ~lo0062;
  assign new_n3929_ = new_n3608_ & new_n3758_;
  assign new_n3930_ = new_n3759_ & new_n3929_;
  assign new_n3931_ = new_n3928_ & new_n3930_;
  assign new_n3932_ = lo0091 & new_n3553_;
  assign new_n3933_ = ~lo0036 & new_n3548_;
  assign new_n3934_ = new_n3748_ & new_n3932_;
  assign new_n3935_ = new_n3547_ & new_n3934_;
  assign new_n3936_ = new_n3933_ & new_n3935_;
  assign new_n3937_ = lo0072 & ~lo0103;
  assign new_n3938_ = new_n3764_ & new_n3937_;
  assign new_n3939_ = new_n3748_ & new_n3813_;
  assign new_n3940_ = new_n3938_ & new_n3939_;
  assign new_n3941_ = ~new_n3936_ & ~new_n3940_;
  assign new_n3942_ = ~new_n3927_ & ~new_n3931_;
  assign new_n3943_ = new_n3941_ & new_n3942_;
  assign new_n3944_ = new_n3924_ & new_n3943_;
  assign new_n3945_ = new_n3608_ & new_n3634_;
  assign new_n3946_ = new_n3580_ & new_n3945_;
  assign new_n3947_ = lo0055 & new_n3946_;
  assign new_n3948_ = new_n3758_ & new_n3947_;
  assign new_n3949_ = ~lo0045 & new_n3573_;
  assign new_n3950_ = new_n3580_ & new_n3949_;
  assign new_n3951_ = lo0053 & new_n3950_;
  assign new_n3952_ = new_n3608_ & new_n3951_;
  assign new_n3953_ = new_n3874_ & new_n3952_;
  assign new_n3954_ = ~new_n3948_ & ~new_n3953_;
  assign new_n3955_ = new_n3557_ & new_n3569_;
  assign new_n3956_ = new_n3716_ & new_n3955_;
  assign new_n3957_ = ~lo0084 & new_n3956_;
  assign new_n3958_ = lo0051 & new_n3957_;
  assign new_n3959_ = new_n3722_ & new_n3958_;
  assign new_n3960_ = lo0109 & new_n3791_;
  assign new_n3961_ = ~lo0069 & new_n3960_;
  assign new_n3962_ = new_n3722_ & new_n3961_;
  assign new_n3963_ = ~new_n3959_ & ~new_n3962_;
  assign new_n3964_ = ~lo0054 & lo0106;
  assign new_n3965_ = new_n3608_ & new_n3964_;
  assign new_n3966_ = new_n3873_ & new_n3965_;
  assign new_n3967_ = new_n3572_ & new_n3709_;
  assign new_n3968_ = new_n3580_ & new_n3967_;
  assign new_n3969_ = new_n3966_ & new_n3968_;
  assign new_n3970_ = new_n3963_ & ~new_n3969_;
  assign new_n3971_ = new_n3590_ & new_n3808_;
  assign new_n3972_ = ~lo0095 & lo0097;
  assign new_n3973_ = new_n3533_ & new_n3971_;
  assign new_n3974_ = new_n3972_ & new_n3973_;
  assign new_n3975_ = new_n3563_ & new_n3565_;
  assign new_n3976_ = ~lo0086 & new_n3569_;
  assign new_n3977_ = new_n3722_ & new_n3975_;
  assign new_n3978_ = new_n3976_ & new_n3977_;
  assign new_n3979_ = lo0077 & new_n3978_;
  assign new_n3980_ = ~new_n3974_ & ~new_n3979_;
  assign new_n3981_ = lo0111 & new_n3553_;
  assign new_n3982_ = new_n3764_ & new_n3981_;
  assign new_n3983_ = ~lo0087 & new_n3982_;
  assign new_n3984_ = new_n3542_ & new_n3983_;
  assign new_n3985_ = new_n3748_ & new_n3984_;
  assign new_n3986_ = ~lo0058 & new_n3550_;
  assign new_n3987_ = lo0098 & new_n3551_;
  assign new_n3988_ = new_n3751_ & new_n3986_;
  assign new_n3989_ = new_n3987_ & new_n3988_;
  assign new_n3990_ = ~new_n3985_ & ~new_n3989_;
  assign new_n3991_ = new_n3980_ & new_n3990_;
  assign new_n3992_ = ~lo0110 & new_n3544_;
  assign new_n3993_ = new_n3829_ & new_n3992_;
  assign new_n3994_ = new_n3553_ & new_n3993_;
  assign new_n3995_ = lo0047 & new_n3994_;
  assign new_n3996_ = new_n3748_ & new_n3995_;
  assign new_n3997_ = ~lo0047 & new_n3553_;
  assign new_n3998_ = new_n3829_ & new_n3997_;
  assign new_n3999_ = lo0110 & new_n3998_;
  assign new_n4000_ = new_n3544_ & new_n3999_;
  assign new_n4001_ = new_n3748_ & new_n4000_;
  assign new_n4002_ = lo0108 & new_n3596_;
  assign new_n4003_ = ~lo0089 & new_n4002_;
  assign new_n4004_ = new_n3530_ & new_n4003_;
  assign new_n4005_ = ~lo0093 & new_n3859_;
  assign new_n4006_ = lo0092 & new_n4005_;
  assign new_n4007_ = new_n3748_ & new_n4006_;
  assign new_n4008_ = ~new_n4004_ & ~new_n4007_;
  assign new_n4009_ = ~new_n4001_ & new_n4008_;
  assign new_n4010_ = new_n3970_ & new_n3991_;
  assign new_n4011_ = ~new_n3996_ & new_n4010_;
  assign new_n4012_ = new_n4009_ & new_n4011_;
  assign new_n4013_ = new_n3954_ & new_n4012_;
  assign new_n4014_ = ~lo0068 & new_n3569_;
  assign new_n4015_ = new_n3741_ & new_n4014_;
  assign new_n4016_ = new_n3560_ & new_n4015_;
  assign new_n4017_ = lo0102 & new_n4016_;
  assign new_n4018_ = new_n3909_ & new_n4017_;
  assign new_n4019_ = lo0095 & new_n3973_;
  assign new_n4020_ = ~lo0097 & new_n4019_;
  assign new_n4021_ = lo0032 & ~lo0038;
  assign new_n4022_ = new_n3606_ & new_n3697_;
  assign new_n4023_ = new_n4021_ & new_n4022_;
  assign new_n4024_ = ~new_n4020_ & ~new_n4023_;
  assign new_n4025_ = ~new_n4018_ & new_n4024_;
  assign new_n4026_ = new_n4013_ & new_n4025_;
  assign new_n4027_ = new_n3944_ & new_n4026_;
  assign new_n4028_ = new_n3729_ & new_n3883_;
  assign new_n4029_ = new_n4027_ & new_n4028_;
  assign new_n4030_ = ~lo0105 & lo0228;
  assign li0025 = ~new_n4029_ & ~new_n4030_;
  assign new_n4032_ = ~new_n3525_ & ~li0025;
  assign new_n4033_ = ~new_n3522_ & new_n4032_;
  assign new_n4034_ = new_n3740_ & ~new_n4020_;
  assign new_n4035_ = ~new_n3746_ & new_n4034_;
  assign new_n4036_ = ~new_n3777_ & ~new_n3794_;
  assign new_n4037_ = ~new_n3769_ & new_n4036_;
  assign new_n4038_ = ~lo0055 & new_n3580_;
  assign new_n4039_ = lo0057 & new_n3520_;
  assign new_n4040_ = new_n3929_ & new_n4038_;
  assign new_n4041_ = new_n4039_ & new_n4040_;
  assign new_n4042_ = new_n4037_ & ~new_n4041_;
  assign new_n4043_ = ~new_n3763_ & ~new_n3773_;
  assign new_n4044_ = new_n4042_ & new_n4043_;
  assign new_n4045_ = new_n3917_ & new_n4044_;
  assign new_n4046_ = ~new_n3780_ & new_n4045_;
  assign new_n4047_ = lo0137 & ~new_n4046_;
  assign new_n4048_ = ~lo0094 & new_n3527_;
  assign new_n4049_ = lo0075 & new_n4048_;
  assign new_n4050_ = new_n3704_ & new_n4049_;
  assign new_n4051_ = lo0198 & ~new_n3636_;
  assign new_n4052_ = ~lo0198 & lo0210;
  assign new_n4053_ = ~new_n4051_ & ~new_n4052_;
  assign new_n4054_ = ~new_n3655_ & new_n4053_;
  assign new_n4055_ = ~lo0137 & ~new_n4054_;
  assign new_n4056_ = new_n4050_ & ~new_n4055_;
  assign new_n4057_ = lo0137 & new_n3799_;
  assign new_n4058_ = ~new_n4056_ & ~new_n4057_;
  assign new_n4059_ = ~new_n4047_ & new_n4058_;
  assign new_n4060_ = ~new_n3786_ & new_n4059_;
  assign new_n4061_ = lo0137 & ~new_n4035_;
  assign new_n4062_ = new_n4060_ & ~new_n4061_;
  assign new_n4063_ = new_n3613_ & ~new_n3753_;
  assign new_n4064_ = ~new_n3828_ & ~new_n3862_;
  assign new_n4065_ = ~new_n3834_ & new_n4064_;
  assign new_n4066_ = new_n3590_ & new_n3809_;
  assign new_n4067_ = ~lo0096 & new_n4066_;
  assign new_n4068_ = lo0074 & new_n4067_;
  assign new_n4069_ = ~new_n3618_ & ~new_n4068_;
  assign new_n4070_ = ~new_n3820_ & ~new_n3879_;
  assign new_n4071_ = new_n4069_ & new_n4070_;
  assign new_n4072_ = ~new_n3870_ & new_n4065_;
  assign new_n4073_ = new_n4071_ & new_n4072_;
  assign new_n4074_ = lo0137 & ~new_n4073_;
  assign new_n4075_ = li0683 & ~new_n4055_;
  assign new_n4076_ = lo0137 & ~li0683;
  assign new_n4077_ = ~new_n4075_ & ~new_n4076_;
  assign new_n4078_ = ~lo0137 & lo0841;
  assign new_n4079_ = lo0137 & new_n4077_;
  assign new_n4080_ = ~new_n4078_ & ~new_n4079_;
  assign new_n4081_ = lo0332 & new_n3804_;
  assign new_n4082_ = lo0137 & new_n3857_;
  assign new_n4083_ = ~new_n4081_ & ~new_n4082_;
  assign new_n4084_ = new_n3810_ & new_n4080_;
  assign new_n4085_ = new_n4083_ & ~new_n4084_;
  assign new_n4086_ = lo0059 & ~lo0060;
  assign new_n4087_ = new_n3733_ & new_n4086_;
  assign new_n4088_ = new_n3783_ & new_n4087_;
  assign new_n4089_ = ~new_n3815_ & ~new_n4088_;
  assign new_n4090_ = lo0137 & ~new_n4089_;
  assign new_n4091_ = lo0841 & ~new_n4053_;
  assign new_n4092_ = lo0225 & new_n4091_;
  assign new_n4093_ = lo0225 & new_n3867_;
  assign new_n4094_ = new_n4023_ & new_n4092_;
  assign new_n4095_ = ~new_n4093_ & ~new_n4094_;
  assign new_n4096_ = lo0841 & new_n4053_;
  assign new_n4097_ = ~new_n4091_ & ~new_n4096_;
  assign new_n4098_ = new_n4023_ & new_n4097_;
  assign new_n4099_ = lo0225 & new_n4098_;
  assign new_n4100_ = lo0137 & ~new_n3847_;
  assign new_n4101_ = ~new_n4099_ & ~new_n4100_;
  assign new_n4102_ = new_n4095_ & new_n4101_;
  assign new_n4103_ = ~new_n4074_ & new_n4085_;
  assign new_n4104_ = ~new_n4090_ & new_n4103_;
  assign new_n4105_ = new_n4102_ & new_n4104_;
  assign new_n4106_ = lo0137 & ~new_n4063_;
  assign new_n4107_ = new_n4105_ & ~new_n4106_;
  assign new_n4108_ = ~new_n3723_ & ~new_n3936_;
  assign new_n4109_ = ~new_n3725_ & new_n4108_;
  assign new_n4110_ = ~new_n3940_ & new_n4109_;
  assign new_n4111_ = lo0137 & new_n3714_;
  assign new_n4112_ = new_n3699_ & ~new_n4055_;
  assign new_n4113_ = ~new_n4111_ & ~new_n4112_;
  assign new_n4114_ = lo0137 & ~new_n4110_;
  assign new_n4115_ = new_n4113_ & ~new_n4114_;
  assign new_n4116_ = ~new_n3922_ & ~new_n4018_;
  assign new_n4117_ = ~new_n3625_ & ~new_n3927_;
  assign new_n4118_ = new_n4116_ & new_n4117_;
  assign new_n4119_ = ~new_n3705_ & ~new_n3931_;
  assign new_n4120_ = new_n4118_ & new_n4119_;
  assign new_n4121_ = lo0137 & ~new_n4120_;
  assign new_n4122_ = new_n4062_ & new_n4107_;
  assign new_n4123_ = new_n4115_ & new_n4122_;
  assign new_n4124_ = ~new_n4121_ & new_n4123_;
  assign new_n4125_ = ~new_n3996_ & ~new_n4001_;
  assign new_n4126_ = ~new_n3959_ & ~new_n3979_;
  assign new_n4127_ = new_n4125_ & new_n4126_;
  assign new_n4128_ = new_n3990_ & new_n4127_;
  assign new_n4129_ = lo0137 & ~new_n4128_;
  assign new_n4130_ = lo0054 & ~lo0106;
  assign new_n4131_ = new_n3608_ & new_n4130_;
  assign new_n4132_ = new_n3873_ & new_n4131_;
  assign new_n4133_ = new_n3968_ & new_n4132_;
  assign new_n4134_ = new_n4008_ & ~new_n4133_;
  assign new_n4135_ = li0683 & ~li0583;
  assign new_n4136_ = ~new_n4055_ & new_n4135_;
  assign new_n4137_ = lo0137 & ~new_n4135_;
  assign new_n4138_ = ~new_n4136_ & ~new_n4137_;
  assign new_n4139_ = new_n3974_ & ~new_n4138_;
  assign new_n4140_ = lo0137 & ~new_n4134_;
  assign new_n4141_ = ~new_n4139_ & ~new_n4140_;
  assign new_n4142_ = ~new_n3962_ & ~new_n3969_;
  assign new_n4143_ = lo0137 & ~new_n4142_;
  assign new_n4144_ = new_n3954_ & ~new_n4129_;
  assign new_n4145_ = new_n4141_ & new_n4144_;
  assign new_n4146_ = ~new_n4143_ & new_n4145_;
  assign li0225 = ~new_n4124_ | ~new_n4146_;
  assign new_n4148_ = lo0095 & ~lo0479;
  assign new_n4149_ = ~lo0040 & ~lo0102;
  assign new_n4150_ = new_n3559_ & new_n4149_;
  assign new_n4151_ = ~lo0055 & ~lo0059;
  assign new_n4152_ = ~lo0062 & new_n4151_;
  assign new_n4153_ = ~lo0060 & new_n3581_;
  assign new_n4154_ = ~lo0056 & ~lo0057;
  assign new_n4155_ = new_n4152_ & new_n4153_;
  assign new_n4156_ = new_n3574_ & new_n4155_;
  assign new_n4157_ = new_n4154_ & new_n4156_;
  assign new_n4158_ = ~lo0032 & ~lo0050;
  assign new_n4159_ = new_n4157_ & new_n4158_;
  assign new_n4160_ = new_n4150_ & new_n4159_;
  assign new_n4161_ = ~lo0100 & new_n4160_;
  assign new_n4162_ = ~lo0038 & new_n4161_;
  assign new_n4163_ = ~lo0069 & ~lo0086;
  assign new_n4164_ = ~lo0077 & ~lo0109;
  assign new_n4165_ = new_n4163_ & new_n4164_;
  assign new_n4166_ = ~lo0087 & ~lo0103;
  assign new_n4167_ = new_n4165_ & new_n4166_;
  assign new_n4168_ = ~lo0104 & ~lo0110;
  assign new_n4169_ = ~lo0088 & new_n4168_;
  assign new_n4170_ = ~lo0047 & new_n4169_;
  assign new_n4171_ = ~lo0072 & ~lo0111;
  assign new_n4172_ = new_n4167_ & new_n4170_;
  assign new_n4173_ = new_n3550_ & new_n4172_;
  assign new_n4174_ = new_n4171_ & new_n4173_;
  assign new_n4175_ = ~lo0071 & ~lo0085;
  assign new_n4176_ = ~lo0067 & ~lo0083;
  assign new_n4177_ = new_n4175_ & new_n4176_;
  assign new_n4178_ = ~lo0068 & ~lo0081;
  assign new_n4179_ = new_n4177_ & new_n4178_;
  assign new_n4180_ = ~lo0065 & new_n4179_;
  assign new_n4181_ = ~li0893 & new_n4180_;
  assign new_n4182_ = ~lo0075 & ~lo0076;
  assign new_n4183_ = ~lo0058 & ~lo0092;
  assign new_n4184_ = ~lo0093 & ~lo0098;
  assign new_n4185_ = new_n4183_ & new_n4184_;
  assign new_n4186_ = ~lo0074 & ~lo0097;
  assign new_n4187_ = new_n4182_ & new_n4185_;
  assign new_n4188_ = new_n4186_ & new_n4187_;
  assign new_n4189_ = ~lo0089 & ~lo0095;
  assign new_n4190_ = ~lo0048 & new_n4189_;
  assign new_n4191_ = lo0096 & new_n4190_;
  assign new_n4192_ = new_n4188_ & new_n4191_;
  assign new_n4193_ = ~lo0039 & ~lo0108;
  assign new_n4194_ = new_n3526_ & new_n4193_;
  assign new_n4195_ = ~lo0049 & ~lo0094;
  assign new_n4196_ = new_n4192_ & new_n4194_;
  assign new_n4197_ = ~lo0095 & new_n4196_;
  assign new_n4198_ = new_n4195_ & new_n4197_;
  assign new_n4199_ = new_n4162_ & new_n4174_;
  assign new_n4200_ = new_n4181_ & new_n4199_;
  assign new_n4201_ = new_n4198_ & new_n4200_;
  assign new_n4202_ = ~new_n4148_ & ~new_n4201_;
  assign new_n4203_ = lo0234 & new_n4202_;
  assign new_n4204_ = ~lo0234 & li0225;
  assign new_n4205_ = ~new_n4203_ & ~new_n4204_;
  assign new_n4206_ = ~new_n3522_ & ~li0025;
  assign new_n4207_ = ~new_n4205_ & ~new_n4206_;
  assign new_n4208_ = ~new_n4033_ & ~new_n4207_;
  assign new_n4209_ = lo0224 & new_n3522_;
  assign new_n4210_ = lo0216 & ~new_n3522_;
  assign new_n4211_ = ~new_n4209_ & ~new_n4210_;
  assign new_n4212_ = lo0222 & ~new_n3522_;
  assign new_n4213_ = lo0221 & ~lo0222;
  assign new_n4214_ = ~new_n4212_ & ~new_n4213_;
  assign new_n4215_ = lo0215 & ~new_n3522_;
  assign new_n4216_ = lo0223 & new_n3522_;
  assign new_n4217_ = ~new_n4215_ & ~new_n4216_;
  assign new_n4218_ = new_n4214_ & new_n4217_;
  assign new_n4219_ = new_n4211_ & new_n4218_;
  assign new_n4220_ = ~new_n4208_ & new_n4219_;
  assign new_n4221_ = ~new_n4214_ & new_n4217_;
  assign new_n4222_ = lo0833 & new_n4221_;
  assign new_n4223_ = new_n4211_ & new_n4222_;
  assign new_n4224_ = lo0929 & new_n4223_;
  assign new_n4225_ = pi055 & ~new_n4223_;
  assign new_n4226_ = ~new_n4224_ & ~new_n4225_;
  assign new_n4227_ = ~new_n4218_ & ~new_n4226_;
  assign new_n4228_ = ~new_n4211_ & new_n4218_;
  assign new_n4229_ = lo0265 & new_n4228_;
  assign new_n4230_ = ~new_n4220_ & ~new_n4227_;
  assign new_n4231_ = ~lo0332 & new_n4230_;
  assign li0000 = new_n4229_ | ~new_n4231_;
  assign new_n4233_ = lo0176 & ~new_n3522_;
  assign new_n4234_ = lo0154 & ~lo0176;
  assign new_n4235_ = ~new_n4233_ & ~new_n4234_;
  assign new_n4236_ = new_n4206_ & new_n4235_;
  assign new_n4237_ = lo0239 & ~new_n4202_;
  assign new_n4238_ = ~new_n4206_ & ~new_n4237_;
  assign new_n4239_ = new_n4219_ & ~new_n4236_;
  assign new_n4240_ = ~new_n4238_ & new_n4239_;
  assign new_n4241_ = lo0276 & new_n4228_;
  assign new_n4242_ = lo0939 & new_n4223_;
  assign new_n4243_ = pi057 & ~new_n4223_;
  assign new_n4244_ = ~new_n4242_ & ~new_n4243_;
  assign new_n4245_ = ~new_n4218_ & ~new_n4244_;
  assign new_n4246_ = ~new_n4240_ & ~new_n4241_;
  assign li0001 = new_n4245_ | ~new_n4246_;
  assign new_n4248_ = ~lo0173 & ~new_n3522_;
  assign new_n4249_ = ~lo0151 & lo0173;
  assign new_n4250_ = ~new_n4248_ & ~new_n4249_;
  assign new_n4251_ = new_n4206_ & ~new_n4250_;
  assign new_n4252_ = lo0235 & ~new_n4202_;
  assign new_n4253_ = ~new_n4206_ & ~new_n4252_;
  assign new_n4254_ = new_n4219_ & ~new_n4251_;
  assign new_n4255_ = ~new_n4253_ & new_n4254_;
  assign new_n4256_ = lo0274 & new_n4228_;
  assign new_n4257_ = lo0927 & new_n4223_;
  assign new_n4258_ = pi056 & ~new_n4223_;
  assign new_n4259_ = ~new_n4257_ & ~new_n4258_;
  assign new_n4260_ = ~new_n4218_ & ~new_n4259_;
  assign new_n4261_ = ~new_n4255_ & ~new_n4256_;
  assign li0002 = new_n4260_ | ~new_n4261_;
  assign new_n4263_ = lo0238 & new_n4202_;
  assign new_n4264_ = ~lo0238 & lo0284;
  assign new_n4265_ = ~new_n4263_ & ~new_n4264_;
  assign new_n4266_ = ~new_n3653_ & ~new_n4206_;
  assign new_n4267_ = new_n3653_ & ~new_n4265_;
  assign new_n4268_ = ~new_n4266_ & ~new_n4267_;
  assign new_n4269_ = new_n4219_ & ~new_n4268_;
  assign new_n4270_ = lo0264 & new_n4228_;
  assign new_n4271_ = ~new_n4269_ & ~new_n4270_;
  assign new_n4272_ = lo0944 & new_n4223_;
  assign new_n4273_ = pi054 & ~new_n4223_;
  assign new_n4274_ = ~new_n4272_ & ~new_n4273_;
  assign new_n4275_ = ~new_n4218_ & ~new_n4274_;
  assign li0003 = ~new_n4271_ | new_n4275_;
  assign new_n4277_ = lo0172 & ~new_n3522_;
  assign new_n4278_ = lo0193 & new_n3522_;
  assign new_n4279_ = ~new_n4277_ & ~new_n4278_;
  assign new_n4280_ = lo0249 & new_n4202_;
  assign new_n4281_ = ~lo0249 & lo0262;
  assign new_n4282_ = ~new_n4280_ & ~new_n4281_;
  assign new_n4283_ = ~new_n4206_ & ~new_n4279_;
  assign new_n4284_ = new_n4279_ & ~new_n4282_;
  assign new_n4285_ = ~new_n4283_ & ~new_n4284_;
  assign new_n4286_ = new_n4219_ & ~new_n4285_;
  assign new_n4287_ = lo0277 & new_n4228_;
  assign new_n4288_ = ~new_n4286_ & ~new_n4287_;
  assign new_n4289_ = lo0932 & new_n4223_;
  assign new_n4290_ = pi053 & ~new_n4223_;
  assign new_n4291_ = ~new_n4289_ & ~new_n4290_;
  assign new_n4292_ = ~new_n4218_ & ~new_n4291_;
  assign li0004 = ~new_n4288_ | new_n4292_;
  assign new_n4294_ = lo0171 & ~new_n3522_;
  assign new_n4295_ = lo0192 & new_n3522_;
  assign new_n4296_ = ~new_n4294_ & ~new_n4295_;
  assign new_n4297_ = lo0241 & new_n4202_;
  assign new_n4298_ = ~lo0241 & lo0861;
  assign new_n4299_ = ~new_n4297_ & ~new_n4298_;
  assign new_n4300_ = ~new_n4206_ & ~new_n4296_;
  assign new_n4301_ = new_n4296_ & ~new_n4299_;
  assign new_n4302_ = ~new_n4300_ & ~new_n4301_;
  assign new_n4303_ = new_n4219_ & ~new_n4302_;
  assign new_n4304_ = lo0270 & new_n4228_;
  assign new_n4305_ = ~new_n4303_ & ~new_n4304_;
  assign new_n4306_ = lo0935 & new_n4223_;
  assign new_n4307_ = pi052 & ~new_n4223_;
  assign new_n4308_ = ~new_n4306_ & ~new_n4307_;
  assign new_n4309_ = ~new_n4218_ & ~new_n4308_;
  assign li0005 = ~new_n4305_ | new_n4309_;
  assign new_n4311_ = lo0170 & ~new_n3522_;
  assign new_n4312_ = lo0194 & new_n3522_;
  assign new_n4313_ = ~new_n4311_ & ~new_n4312_;
  assign new_n4314_ = lo0248 & new_n4202_;
  assign new_n4315_ = ~lo0248 & lo0869;
  assign new_n4316_ = ~new_n4314_ & ~new_n4315_;
  assign new_n4317_ = ~new_n4206_ & ~new_n4313_;
  assign new_n4318_ = new_n4313_ & ~new_n4316_;
  assign new_n4319_ = ~new_n4317_ & ~new_n4318_;
  assign new_n4320_ = new_n4219_ & ~new_n4319_;
  assign new_n4321_ = lo0282 & new_n4228_;
  assign new_n4322_ = ~new_n4320_ & ~new_n4321_;
  assign new_n4323_ = lo0921 & new_n4223_;
  assign new_n4324_ = pi051 & ~new_n4223_;
  assign new_n4325_ = ~new_n4323_ & ~new_n4324_;
  assign new_n4326_ = ~new_n4218_ & ~new_n4325_;
  assign li0006 = ~new_n4322_ | new_n4326_;
  assign new_n4328_ = lo0141 & new_n3522_;
  assign new_n4329_ = lo0148 & ~new_n3522_;
  assign new_n4330_ = ~new_n4328_ & ~new_n4329_;
  assign new_n4331_ = lo0247 & new_n4202_;
  assign new_n4332_ = ~lo0247 & lo0862;
  assign new_n4333_ = ~new_n4331_ & ~new_n4332_;
  assign new_n4334_ = ~new_n4206_ & ~new_n4330_;
  assign new_n4335_ = new_n4330_ & ~new_n4333_;
  assign new_n4336_ = ~new_n4334_ & ~new_n4335_;
  assign new_n4337_ = new_n4219_ & ~new_n4336_;
  assign new_n4338_ = lo0281 & new_n4228_;
  assign new_n4339_ = ~new_n4337_ & ~new_n4338_;
  assign new_n4340_ = lo0920 & new_n4223_;
  assign new_n4341_ = pi050 & ~new_n4223_;
  assign new_n4342_ = ~new_n4340_ & ~new_n4341_;
  assign new_n4343_ = ~new_n4218_ & ~new_n4342_;
  assign li0007 = ~new_n4339_ | new_n4343_;
  assign new_n4345_ = lo0191 & new_n3522_;
  assign new_n4346_ = lo0169 & ~new_n3522_;
  assign new_n4347_ = ~new_n4345_ & ~new_n4346_;
  assign new_n4348_ = lo0246 & new_n4202_;
  assign new_n4349_ = ~lo0246 & lo0877;
  assign new_n4350_ = ~new_n4348_ & ~new_n4349_;
  assign new_n4351_ = ~new_n4206_ & ~new_n4347_;
  assign new_n4352_ = new_n4347_ & ~new_n4350_;
  assign new_n4353_ = ~new_n4351_ & ~new_n4352_;
  assign new_n4354_ = new_n4219_ & ~new_n4353_;
  assign new_n4355_ = lo0269 & new_n4228_;
  assign new_n4356_ = ~new_n4354_ & ~new_n4355_;
  assign new_n4357_ = lo0940 & new_n4223_;
  assign new_n4358_ = pi049 & ~new_n4223_;
  assign new_n4359_ = ~new_n4357_ & ~new_n4358_;
  assign new_n4360_ = ~new_n4218_ & ~new_n4359_;
  assign li0008 = ~new_n4356_ | new_n4360_;
  assign new_n4362_ = lo0168 & ~new_n3522_;
  assign new_n4363_ = lo0190 & new_n3522_;
  assign new_n4364_ = ~new_n4362_ & ~new_n4363_;
  assign new_n4365_ = lo0240 & new_n4202_;
  assign new_n4366_ = ~lo0240 & lo0878;
  assign new_n4367_ = ~new_n4365_ & ~new_n4366_;
  assign new_n4368_ = ~new_n4206_ & ~new_n4364_;
  assign new_n4369_ = new_n4364_ & ~new_n4367_;
  assign new_n4370_ = ~new_n4368_ & ~new_n4369_;
  assign new_n4371_ = new_n4219_ & ~new_n4370_;
  assign new_n4372_ = lo0280 & new_n4228_;
  assign new_n4373_ = ~new_n4371_ & ~new_n4372_;
  assign new_n4374_ = lo0933 & new_n4223_;
  assign new_n4375_ = pi048 & ~new_n4223_;
  assign new_n4376_ = ~new_n4374_ & ~new_n4375_;
  assign new_n4377_ = ~new_n4218_ & ~new_n4376_;
  assign li0009 = ~new_n4373_ | new_n4377_;
  assign new_n4379_ = lo0245 & new_n4202_;
  assign new_n4380_ = ~lo0245 & lo0875;
  assign new_n4381_ = ~new_n4379_ & ~new_n4380_;
  assign new_n4382_ = ~new_n3645_ & ~new_n4206_;
  assign new_n4383_ = new_n3645_ & ~new_n4381_;
  assign new_n4384_ = ~new_n4382_ & ~new_n4383_;
  assign new_n4385_ = new_n4219_ & ~new_n4384_;
  assign new_n4386_ = lo0266 & new_n4228_;
  assign new_n4387_ = ~new_n4385_ & ~new_n4386_;
  assign new_n4388_ = lo0928 & new_n4223_;
  assign new_n4389_ = pi047 & ~new_n4223_;
  assign new_n4390_ = ~new_n4388_ & ~new_n4389_;
  assign new_n4391_ = ~new_n4218_ & ~new_n4390_;
  assign li0010 = ~new_n4387_ | new_n4391_;
  assign new_n4393_ = lo0244 & new_n4202_;
  assign new_n4394_ = ~lo0244 & lo0879;
  assign new_n4395_ = ~new_n4393_ & ~new_n4394_;
  assign new_n4396_ = ~new_n3639_ & ~new_n4206_;
  assign new_n4397_ = new_n3639_ & ~new_n4395_;
  assign new_n4398_ = ~new_n4396_ & ~new_n4397_;
  assign new_n4399_ = new_n4219_ & ~new_n4398_;
  assign new_n4400_ = lo0279 & new_n4228_;
  assign new_n4401_ = ~new_n4399_ & ~new_n4400_;
  assign new_n4402_ = lo0938 & new_n4223_;
  assign new_n4403_ = pi046 & ~new_n4223_;
  assign new_n4404_ = ~new_n4402_ & ~new_n4403_;
  assign new_n4405_ = ~new_n4218_ & ~new_n4404_;
  assign li0011 = ~new_n4401_ | new_n4405_;
  assign new_n4407_ = lo0242 & new_n4202_;
  assign new_n4408_ = ~lo0242 & lo0846;
  assign new_n4409_ = ~new_n4407_ & ~new_n4408_;
  assign new_n4410_ = ~new_n3633_ & ~new_n4206_;
  assign new_n4411_ = new_n3633_ & ~new_n4409_;
  assign new_n4412_ = ~new_n4410_ & ~new_n4411_;
  assign new_n4413_ = new_n4219_ & ~new_n4412_;
  assign new_n4414_ = lo0278 & new_n4228_;
  assign new_n4415_ = ~new_n4413_ & ~new_n4414_;
  assign new_n4416_ = lo0930 & new_n4223_;
  assign new_n4417_ = pi045 & ~new_n4223_;
  assign new_n4418_ = ~new_n4416_ & ~new_n4417_;
  assign new_n4419_ = ~new_n4218_ & ~new_n4418_;
  assign li0012 = ~new_n4415_ | new_n4419_;
  assign new_n4421_ = lo0835 & lo0984;
  assign new_n4422_ = ~lo0979 & ~new_n4421_;
  assign new_n4423_ = ~lo0252 & lo0995;
  assign new_n4424_ = new_n4422_ & ~new_n4423_;
  assign new_n4425_ = ~new_n4219_ & ~new_n4228_;
  assign new_n4426_ = new_n4211_ & new_n4217_;
  assign new_n4427_ = ~new_n4214_ & new_n4426_;
  assign new_n4428_ = ~new_n4211_ & new_n4221_;
  assign new_n4429_ = lo0969 & new_n3636_;
  assign new_n4430_ = lo0963 & ~new_n3522_;
  assign new_n4431_ = ~new_n4429_ & ~new_n4430_;
  assign new_n4432_ = lo0967 & new_n3636_;
  assign new_n4433_ = lo0970 & ~new_n3522_;
  assign new_n4434_ = ~new_n4432_ & ~new_n4433_;
  assign new_n4435_ = lo0977 & new_n3522_;
  assign new_n4436_ = lo0960 & ~new_n3522_;
  assign new_n4437_ = ~new_n4435_ & ~new_n4436_;
  assign new_n4438_ = lo0961 & new_n3522_;
  assign new_n4439_ = lo0972 & ~new_n3636_;
  assign new_n4440_ = ~new_n4438_ & ~new_n4439_;
  assign new_n4441_ = new_n4431_ & new_n4434_;
  assign new_n4442_ = new_n4437_ & new_n4441_;
  assign new_n4443_ = new_n4440_ & new_n4442_;
  assign new_n4444_ = new_n3641_ & ~new_n4443_;
  assign new_n4445_ = lo0974 & ~new_n3636_;
  assign new_n4446_ = ~lo0974 & lo0978;
  assign new_n4447_ = ~new_n4445_ & ~new_n4446_;
  assign new_n4448_ = lo0971 & ~new_n3636_;
  assign new_n4449_ = ~lo0971 & lo0975;
  assign new_n4450_ = ~new_n4448_ & ~new_n4449_;
  assign new_n4451_ = new_n4447_ & new_n4450_;
  assign new_n4452_ = ~lo0614 & ~lo0642;
  assign new_n4453_ = ~lo0616 & new_n4452_;
  assign new_n4454_ = lo0603 & new_n4453_;
  assign new_n4455_ = lo0587 & new_n3522_;
  assign new_n4456_ = lo0947 & ~new_n3636_;
  assign new_n4457_ = ~new_n4455_ & ~new_n4456_;
  assign new_n4458_ = new_n3641_ & ~new_n4454_;
  assign new_n4459_ = new_n4454_ & new_n4457_;
  assign new_n4460_ = ~new_n4458_ & ~new_n4459_;
  assign new_n4461_ = lo0602 & ~new_n3522_;
  assign new_n4462_ = ~lo0602 & lo0907;
  assign new_n4463_ = ~new_n4461_ & ~new_n4462_;
  assign new_n4464_ = ~lo0661 & lo0680;
  assign new_n4465_ = ~lo0662 & ~lo0681;
  assign new_n4466_ = new_n4464_ & new_n4465_;
  assign new_n4467_ = ~new_n3641_ & new_n4466_;
  assign new_n4468_ = new_n3641_ & ~new_n4463_;
  assign new_n4469_ = ~new_n4467_ & ~new_n4468_;
  assign new_n4470_ = ~new_n4460_ & new_n4469_;
  assign new_n4471_ = new_n3641_ & ~new_n4451_;
  assign new_n4472_ = new_n4470_ & ~new_n4471_;
  assign new_n4473_ = ~new_n4444_ & new_n4472_;
  assign new_n4474_ = lo0835 & ~li0793;
  assign new_n4475_ = ~new_n4473_ & new_n4474_;
  assign new_n4476_ = ~new_n4135_ & new_n4428_;
  assign new_n4477_ = new_n4475_ & ~new_n4476_;
  assign new_n4478_ = new_n4424_ & new_n4425_;
  assign new_n4479_ = ~new_n4427_ & new_n4478_;
  assign new_n4480_ = new_n4477_ & new_n4479_;
  assign new_n4481_ = new_n3612_ & ~new_n4480_;
  assign new_n4482_ = lo0287 & new_n3612_;
  assign new_n4483_ = ~new_n3589_ & ~new_n4481_;
  assign new_n4484_ = ~new_n4482_ & new_n4483_;
  assign new_n4485_ = ~new_n3828_ & new_n3847_;
  assign new_n4486_ = ~new_n3815_ & new_n4485_;
  assign new_n4487_ = new_n3871_ & new_n4486_;
  assign new_n4488_ = lo0841 & new_n3862_;
  assign new_n4489_ = ~new_n3834_ & ~new_n3857_;
  assign new_n4490_ = ~new_n4488_ & new_n4489_;
  assign new_n4491_ = ~new_n3879_ & new_n4490_;
  assign new_n4492_ = ~new_n3810_ & ~new_n3820_;
  assign new_n4493_ = new_n4069_ & new_n4492_;
  assign new_n4494_ = new_n4491_ & new_n4493_;
  assign new_n4495_ = new_n3755_ & ~new_n4020_;
  assign new_n4496_ = new_n4487_ & new_n4495_;
  assign new_n4497_ = new_n4494_ & new_n4496_;
  assign new_n4498_ = new_n4023_ & new_n4091_;
  assign new_n4499_ = new_n4023_ & ~new_n4096_;
  assign new_n4500_ = ~new_n4498_ & ~new_n4499_;
  assign new_n4501_ = ~new_n3969_ & new_n4045_;
  assign new_n4502_ = ~new_n3962_ & ~new_n3974_;
  assign new_n4503_ = ~new_n3940_ & new_n4119_;
  assign new_n4504_ = ~new_n3668_ & new_n3690_;
  assign new_n4505_ = ~new_n3669_ & new_n4504_;
  assign new_n4506_ = ~new_n3694_ & ~new_n4505_;
  assign new_n4507_ = new_n3699_ & ~new_n4506_;
  assign new_n4508_ = ~new_n3723_ & new_n4503_;
  assign new_n4509_ = new_n3715_ & new_n4508_;
  assign new_n4510_ = ~new_n4507_ & new_n4509_;
  assign new_n4511_ = new_n4118_ & new_n4502_;
  assign new_n4512_ = ~new_n3725_ & new_n4511_;
  assign new_n4513_ = new_n4510_ & new_n4512_;
  assign new_n4514_ = new_n4501_ & new_n4513_;
  assign new_n4515_ = ~new_n4001_ & ~new_n4004_;
  assign new_n4516_ = new_n3990_ & new_n4515_;
  assign new_n4517_ = new_n4514_ & new_n4516_;
  assign new_n4518_ = ~new_n3996_ & new_n4517_;
  assign new_n4519_ = ~new_n3959_ & new_n4518_;
  assign new_n4520_ = new_n4484_ & new_n4497_;
  assign new_n4521_ = new_n4500_ & new_n4520_;
  assign li0013 = ~new_n4519_ | ~new_n4521_;
  assign new_n4523_ = ~lo0479 & new_n4020_;
  assign new_n4524_ = ~lo0287 & ~lo0979;
  assign new_n4525_ = new_n3612_ & new_n4524_;
  assign new_n4526_ = ~new_n4421_ & ~new_n4423_;
  assign new_n4527_ = new_n4525_ & new_n4526_;
  assign new_n4528_ = ~li0683 & ~li0583;
  assign new_n4529_ = new_n4427_ & new_n4528_;
  assign new_n4530_ = ~li0583 & new_n4428_;
  assign new_n4531_ = ~new_n4529_ & ~new_n4530_;
  assign new_n4532_ = new_n4475_ & ~new_n4531_;
  assign new_n4533_ = new_n4527_ & new_n4532_;
  assign new_n4534_ = ~new_n4091_ & new_n4096_;
  assign new_n4535_ = new_n4023_ & new_n4534_;
  assign new_n4536_ = ~new_n4523_ & ~new_n4533_;
  assign new_n4537_ = ~new_n4535_ & new_n4536_;
  assign new_n4538_ = lo0145 & ~new_n3522_;
  assign new_n4539_ = ~lo0145 & lo0197;
  assign new_n4540_ = ~new_n4538_ & ~new_n4539_;
  assign new_n4541_ = ~new_n3630_ & new_n3642_;
  assign new_n4542_ = ~new_n3614_ & new_n4541_;
  assign new_n4543_ = ~new_n3628_ & new_n4542_;
  assign new_n4544_ = new_n4540_ & new_n4543_;
  assign new_n4545_ = lo0181 & ~new_n3522_;
  assign new_n4546_ = lo0159 & ~lo0181;
  assign new_n4547_ = ~new_n4545_ & ~new_n4546_;
  assign new_n4548_ = new_n4543_ & new_n4547_;
  assign new_n4549_ = new_n4544_ & new_n4548_;
  assign new_n4550_ = lo0182 & ~new_n3522_;
  assign new_n4551_ = lo0160 & ~lo0182;
  assign new_n4552_ = ~new_n4550_ & ~new_n4551_;
  assign new_n4553_ = new_n4543_ & new_n4552_;
  assign new_n4554_ = lo0180 & ~new_n3522_;
  assign new_n4555_ = lo0158 & ~lo0180;
  assign new_n4556_ = ~new_n4554_ & ~new_n4555_;
  assign new_n4557_ = new_n4543_ & new_n4556_;
  assign new_n4558_ = new_n4553_ & new_n4557_;
  assign new_n4559_ = new_n4549_ & new_n4558_;
  assign new_n4560_ = new_n3962_ & ~new_n4559_;
  assign new_n4561_ = ~new_n3780_ & ~new_n4050_;
  assign new_n4562_ = ~new_n3799_ & new_n4561_;
  assign new_n4563_ = ~new_n3723_ & new_n4562_;
  assign new_n4564_ = ~new_n3804_ & ~new_n3857_;
  assign new_n4565_ = ~lo0841 & new_n3862_;
  assign new_n4566_ = ~new_n3618_ & ~new_n3870_;
  assign new_n4567_ = ~lo0314 & new_n3815_;
  assign new_n4568_ = ~new_n4088_ & ~new_n4565_;
  assign new_n4569_ = new_n4566_ & new_n4568_;
  assign new_n4570_ = ~new_n4567_ & new_n4569_;
  assign new_n4571_ = new_n4564_ & new_n4570_;
  assign new_n4572_ = ~new_n4068_ & new_n4485_;
  assign new_n4573_ = new_n4563_ & new_n4571_;
  assign new_n4574_ = new_n4572_ & new_n4573_;
  assign new_n4575_ = ~new_n3794_ & ~new_n3914_;
  assign new_n4576_ = ~new_n3898_ & new_n4575_;
  assign new_n4577_ = ~new_n3907_ & new_n4576_;
  assign new_n4578_ = ~new_n3786_ & ~new_n3903_;
  assign new_n4579_ = ~new_n4041_ & new_n4578_;
  assign new_n4580_ = new_n3668_ & ~new_n3688_;
  assign new_n4581_ = ~new_n3689_ & new_n4580_;
  assign new_n4582_ = ~new_n3669_ & ~new_n4581_;
  assign new_n4583_ = new_n3699_ & ~new_n4582_;
  assign new_n4584_ = ~new_n3940_ & ~new_n4583_;
  assign new_n4585_ = ~new_n3936_ & new_n4584_;
  assign new_n4586_ = ~new_n3625_ & new_n4585_;
  assign new_n4587_ = new_n4574_ & new_n4577_;
  assign new_n4588_ = new_n4579_ & new_n4587_;
  assign new_n4589_ = new_n4586_ & new_n4588_;
  assign new_n4590_ = new_n4537_ & ~new_n4560_;
  assign new_n4591_ = new_n4589_ & new_n4590_;
  assign new_n4592_ = ~new_n3746_ & ~new_n4007_;
  assign new_n4593_ = ~new_n3979_ & ~new_n4133_;
  assign new_n4594_ = new_n3954_ & new_n4593_;
  assign new_n4595_ = new_n4591_ & new_n4592_;
  assign li0037 = ~new_n4594_ | ~new_n4595_;
  assign new_n4597_ = ~lo0228 & li0037;
  assign new_n4598_ = lo0030 & lo0228;
  assign new_n4599_ = ~new_n4597_ & ~new_n4598_;
  assign li0014 = new_n4469_ | new_n4599_;
  assign li0015 = ~new_n4460_ | new_n4599_;
  assign new_n4602_ = new_n3641_ & ~new_n4434_;
  assign li0016 = new_n4599_ | ~new_n4602_;
  assign new_n4604_ = new_n3641_ & ~new_n4440_;
  assign li0017 = new_n4599_ | ~new_n4604_;
  assign new_n4606_ = new_n3641_ & ~new_n4437_;
  assign li0018 = new_n4599_ | ~new_n4606_;
  assign new_n4608_ = new_n3641_ & ~new_n4431_;
  assign li0019 = new_n4599_ | ~new_n4608_;
  assign new_n4610_ = new_n3641_ & ~new_n4450_;
  assign li0020 = new_n4599_ | ~new_n4610_;
  assign new_n4612_ = new_n3641_ & ~new_n4447_;
  assign li0021 = new_n4599_ | ~new_n4612_;
  assign new_n4614_ = lo0024 & lo0954;
  assign new_n4615_ = ~lo0954 & li0037;
  assign li0024 = new_n4614_ | new_n4615_;
  assign new_n4617_ = ~lo0228 & lo0252;
  assign new_n4618_ = ~lo0119 & ~new_n4617_;
  assign new_n4619_ = lo0119 & ~lo1050;
  assign new_n4620_ = ~new_n4618_ & ~new_n4619_;
  assign li0026 = lo0468 | ~new_n4620_;
  assign new_n4622_ = lo0119 & ~lo1071;
  assign new_n4623_ = ~new_n4618_ & ~new_n4622_;
  assign li0027 = lo0468 | ~new_n4623_;
  assign new_n4625_ = lo0119 & ~lo1067;
  assign new_n4626_ = ~new_n4618_ & ~new_n4625_;
  assign li0028 = lo0468 | ~new_n4626_;
  assign new_n4628_ = lo0119 & ~lo1035;
  assign new_n4629_ = ~new_n4618_ & ~new_n4628_;
  assign li0029 = lo0468 | ~new_n4629_;
  assign new_n4631_ = lo0024 & new_n3936_;
  assign new_n4632_ = ~lo0122 & ~li0583;
  assign new_n4633_ = new_n4631_ & new_n4632_;
  assign new_n4634_ = li0683 & new_n4633_;
  assign new_n4635_ = ~lo0122 & new_n4135_;
  assign new_n4636_ = new_n3974_ & new_n4635_;
  assign new_n4637_ = lo0841 & new_n3857_;
  assign new_n4638_ = ~new_n3769_ & ~new_n4637_;
  assign new_n4639_ = ~new_n3989_ & new_n4638_;
  assign new_n4640_ = ~new_n3959_ & new_n4639_;
  assign new_n4641_ = ~new_n4488_ & new_n4640_;
  assign new_n4642_ = ~new_n4636_ & new_n4641_;
  assign new_n4643_ = ~new_n4634_ & new_n4642_;
  assign new_n4644_ = ~lo0122 & li0683;
  assign new_n4645_ = ~li0583 & new_n4644_;
  assign new_n4646_ = lo0228 & new_n4645_;
  assign new_n4647_ = ~new_n3650_ & li0901;
  assign new_n4648_ = new_n3699_ & new_n4646_;
  assign new_n4649_ = new_n4647_ & new_n4648_;
  assign new_n4650_ = new_n3810_ & new_n4644_;
  assign new_n4651_ = lo0841 & new_n4650_;
  assign new_n4652_ = ~new_n4649_ & ~new_n4651_;
  assign new_n4653_ = ~lo0287 & new_n3612_;
  assign new_n4654_ = new_n4475_ & new_n4653_;
  assign new_n4655_ = new_n4135_ & new_n4427_;
  assign new_n4656_ = new_n4654_ & new_n4655_;
  assign new_n4657_ = new_n4424_ & new_n4656_;
  assign new_n4658_ = lo0024 & new_n4644_;
  assign new_n4659_ = lo0252 & new_n4658_;
  assign new_n4660_ = new_n4050_ & new_n4659_;
  assign new_n4661_ = ~li0583 & new_n4660_;
  assign new_n4662_ = new_n4647_ & new_n4661_;
  assign new_n4663_ = new_n4643_ & new_n4652_;
  assign new_n4664_ = ~new_n4657_ & new_n4663_;
  assign new_n4665_ = ~new_n4662_ & new_n4664_;
  assign new_n4666_ = pi002 & pi004;
  assign new_n4667_ = ~lo0286 & ~lo0288;
  assign new_n4668_ = ~lo0289 & new_n4667_;
  assign new_n4669_ = ~lo0285 & new_n4668_;
  assign new_n4670_ = new_n4632_ & ~new_n4666_;
  assign new_n4671_ = new_n3678_ & new_n4670_;
  assign new_n4672_ = ~new_n4669_ & new_n4671_;
  assign new_n4673_ = new_n4665_ & ~new_n4672_;
  assign li0122 = ~li0793 & ~new_n4673_;
  assign new_n4675_ = ~pi002 & lo0217;
  assign new_n4676_ = new_n3673_ & new_n4675_;
  assign new_n4677_ = ~li0793 & new_n4676_;
  assign new_n4678_ = ~new_n4673_ & new_n4677_;
  assign new_n4679_ = ~lo0590 & ~lo0592;
  assign new_n4680_ = ~lo0588 & new_n4679_;
  assign new_n4681_ = lo0591 & new_n4680_;
  assign new_n4682_ = lo0588 & ~lo0590;
  assign new_n4683_ = ~lo0591 & ~lo0592;
  assign new_n4684_ = new_n4682_ & new_n4683_;
  assign new_n4685_ = lo0324 & new_n4681_;
  assign new_n4686_ = lo0446 & new_n4684_;
  assign new_n4687_ = ~new_n4685_ & ~new_n4686_;
  assign new_n4688_ = ~lo0588 & ~lo0590;
  assign new_n4689_ = ~lo0591 & new_n4688_;
  assign new_n4690_ = lo0592 & new_n4689_;
  assign new_n4691_ = ~lo0588 & ~lo0591;
  assign new_n4692_ = ~lo0592 & new_n4691_;
  assign new_n4693_ = lo0590 & new_n4692_;
  assign new_n4694_ = lo0339 & new_n4690_;
  assign new_n4695_ = lo0460 & new_n4693_;
  assign new_n4696_ = ~new_n4694_ & ~new_n4695_;
  assign new_n4697_ = new_n4687_ & new_n4696_;
  assign new_n4698_ = lo0456 & new_n4681_;
  assign new_n4699_ = lo0443 & new_n4684_;
  assign new_n4700_ = ~new_n4698_ & ~new_n4699_;
  assign new_n4701_ = lo0337 & new_n4690_;
  assign new_n4702_ = lo0441 & new_n4693_;
  assign new_n4703_ = ~new_n4701_ & ~new_n4702_;
  assign new_n4704_ = new_n4700_ & new_n4703_;
  assign new_n4705_ = lo0390 & new_n4681_;
  assign new_n4706_ = lo0342 & new_n4693_;
  assign new_n4707_ = ~new_n4705_ & ~new_n4706_;
  assign new_n4708_ = lo0414 & new_n4684_;
  assign new_n4709_ = lo0363 & new_n4690_;
  assign new_n4710_ = ~new_n4708_ & ~new_n4709_;
  assign new_n4711_ = new_n4707_ & new_n4710_;
  assign new_n4712_ = new_n4704_ & ~new_n4711_;
  assign new_n4713_ = ~new_n4704_ & new_n4711_;
  assign new_n4714_ = ~new_n4712_ & ~new_n4713_;
  assign new_n4715_ = lo0380 & new_n4690_;
  assign new_n4716_ = lo0355 & new_n4693_;
  assign new_n4717_ = ~new_n4715_ & ~new_n4716_;
  assign new_n4718_ = lo0404 & new_n4681_;
  assign new_n4719_ = lo0429 & new_n4684_;
  assign new_n4720_ = ~new_n4718_ & ~new_n4719_;
  assign new_n4721_ = new_n4717_ & new_n4720_;
  assign new_n4722_ = lo0386 & new_n4690_;
  assign new_n4723_ = lo0361 & new_n4693_;
  assign new_n4724_ = ~new_n4722_ & ~new_n4723_;
  assign new_n4725_ = lo0410 & new_n4681_;
  assign new_n4726_ = lo0434 & new_n4684_;
  assign new_n4727_ = ~new_n4725_ & ~new_n4726_;
  assign new_n4728_ = new_n4724_ & new_n4727_;
  assign new_n4729_ = new_n4721_ & ~new_n4728_;
  assign new_n4730_ = ~new_n4721_ & new_n4728_;
  assign new_n4731_ = ~new_n4729_ & ~new_n4730_;
  assign new_n4732_ = new_n4714_ & ~new_n4731_;
  assign new_n4733_ = ~new_n4714_ & new_n4731_;
  assign new_n4734_ = ~new_n4732_ & ~new_n4733_;
  assign new_n4735_ = lo0319 & new_n4681_;
  assign new_n4736_ = lo0458 & new_n4693_;
  assign new_n4737_ = ~new_n4735_ & ~new_n4736_;
  assign new_n4738_ = lo0444 & new_n4684_;
  assign new_n4739_ = lo0338 & new_n4690_;
  assign new_n4740_ = ~new_n4738_ & ~new_n4739_;
  assign new_n4741_ = new_n4737_ & new_n4740_;
  assign new_n4742_ = lo0411 & new_n4681_;
  assign new_n4743_ = lo0435 & new_n4684_;
  assign new_n4744_ = ~new_n4742_ & ~new_n4743_;
  assign new_n4745_ = lo0387 & new_n4690_;
  assign new_n4746_ = lo0452 & new_n4693_;
  assign new_n4747_ = ~new_n4745_ & ~new_n4746_;
  assign new_n4748_ = new_n4744_ & new_n4747_;
  assign new_n4749_ = new_n4741_ & ~new_n4748_;
  assign new_n4750_ = ~new_n4741_ & new_n4748_;
  assign new_n4751_ = ~new_n4749_ & ~new_n4750_;
  assign new_n4752_ = lo0372 & new_n4690_;
  assign new_n4753_ = lo0320 & new_n4693_;
  assign new_n4754_ = ~new_n4752_ & ~new_n4753_;
  assign new_n4755_ = lo0397 & new_n4681_;
  assign new_n4756_ = lo0422 & new_n4684_;
  assign new_n4757_ = ~new_n4755_ & ~new_n4756_;
  assign new_n4758_ = new_n4754_ & new_n4757_;
  assign new_n4759_ = lo0412 & new_n4681_;
  assign new_n4760_ = lo0388 & new_n4690_;
  assign new_n4761_ = ~new_n4759_ & ~new_n4760_;
  assign new_n4762_ = lo0436 & new_n4684_;
  assign new_n4763_ = lo0455 & new_n4693_;
  assign new_n4764_ = ~new_n4762_ & ~new_n4763_;
  assign new_n4765_ = new_n4761_ & new_n4764_;
  assign new_n4766_ = new_n4758_ & ~new_n4765_;
  assign new_n4767_ = ~new_n4758_ & new_n4765_;
  assign new_n4768_ = ~new_n4766_ & ~new_n4767_;
  assign new_n4769_ = new_n4751_ & ~new_n4768_;
  assign new_n4770_ = ~new_n4751_ & new_n4768_;
  assign new_n4771_ = ~new_n4769_ & ~new_n4770_;
  assign new_n4772_ = new_n4734_ & ~new_n4771_;
  assign new_n4773_ = ~new_n4734_ & new_n4771_;
  assign new_n4774_ = ~new_n4772_ & ~new_n4773_;
  assign new_n4775_ = new_n4697_ & ~new_n4774_;
  assign new_n4776_ = ~new_n4697_ & new_n4774_;
  assign new_n4777_ = ~new_n4775_ & ~new_n4776_;
  assign new_n4778_ = pi107 & ~new_n4777_;
  assign new_n4779_ = lo0384 & new_n4690_;
  assign new_n4780_ = lo0359 & new_n4693_;
  assign new_n4781_ = ~new_n4779_ & ~new_n4780_;
  assign new_n4782_ = lo0408 & new_n4681_;
  assign new_n4783_ = lo0432 & new_n4684_;
  assign new_n4784_ = ~new_n4782_ & ~new_n4783_;
  assign new_n4785_ = new_n4781_ & new_n4784_;
  assign new_n4786_ = lo0396 & new_n4681_;
  assign new_n4787_ = lo0322 & new_n4693_;
  assign new_n4788_ = ~new_n4786_ & ~new_n4787_;
  assign new_n4789_ = lo0421 & new_n4684_;
  assign new_n4790_ = lo0371 & new_n4690_;
  assign new_n4791_ = ~new_n4789_ & ~new_n4790_;
  assign new_n4792_ = new_n4788_ & new_n4791_;
  assign new_n4793_ = lo0349 & new_n4693_;
  assign new_n4794_ = lo0440 & new_n4690_;
  assign new_n4795_ = ~new_n4793_ & ~new_n4794_;
  assign new_n4796_ = lo0329 & new_n4681_;
  assign new_n4797_ = lo0454 & new_n4684_;
  assign new_n4798_ = new_n4795_ & ~new_n4796_;
  assign new_n4799_ = ~new_n4797_ & new_n4798_;
  assign new_n4800_ = new_n4792_ & ~new_n4799_;
  assign new_n4801_ = ~new_n4792_ & new_n4799_;
  assign new_n4802_ = ~new_n4800_ & ~new_n4801_;
  assign new_n4803_ = lo0370 & new_n4690_;
  assign new_n4804_ = lo0347 & new_n4693_;
  assign new_n4805_ = ~new_n4803_ & ~new_n4804_;
  assign new_n4806_ = lo0395 & new_n4681_;
  assign new_n4807_ = lo0420 & new_n4684_;
  assign new_n4808_ = ~new_n4806_ & ~new_n4807_;
  assign new_n4809_ = new_n4805_ & new_n4808_;
  assign new_n4810_ = lo0375 & new_n4690_;
  assign new_n4811_ = lo0316 & new_n4693_;
  assign new_n4812_ = ~new_n4810_ & ~new_n4811_;
  assign new_n4813_ = lo0399 & new_n4681_;
  assign new_n4814_ = lo0424 & new_n4684_;
  assign new_n4815_ = ~new_n4813_ & ~new_n4814_;
  assign new_n4816_ = new_n4812_ & new_n4815_;
  assign new_n4817_ = new_n4809_ & ~new_n4816_;
  assign new_n4818_ = ~new_n4809_ & new_n4816_;
  assign new_n4819_ = ~new_n4817_ & ~new_n4818_;
  assign new_n4820_ = new_n4802_ & ~new_n4819_;
  assign new_n4821_ = ~new_n4802_ & new_n4819_;
  assign new_n4822_ = ~new_n4820_ & ~new_n4821_;
  assign new_n4823_ = lo0374 & new_n4690_;
  assign new_n4824_ = lo0350 & new_n4693_;
  assign new_n4825_ = ~new_n4823_ & ~new_n4824_;
  assign new_n4826_ = lo0400 & new_n4681_;
  assign new_n4827_ = lo0425 & new_n4684_;
  assign new_n4828_ = ~new_n4826_ & ~new_n4827_;
  assign new_n4829_ = new_n4825_ & new_n4828_;
  assign new_n4830_ = lo0369 & new_n4690_;
  assign new_n4831_ = lo0315 & new_n4693_;
  assign new_n4832_ = ~new_n4830_ & ~new_n4831_;
  assign new_n4833_ = lo0394 & new_n4681_;
  assign new_n4834_ = lo0419 & new_n4684_;
  assign new_n4835_ = ~new_n4833_ & ~new_n4834_;
  assign new_n4836_ = new_n4832_ & new_n4835_;
  assign new_n4837_ = new_n4829_ & ~new_n4836_;
  assign new_n4838_ = ~new_n4829_ & new_n4836_;
  assign new_n4839_ = ~new_n4837_ & ~new_n4838_;
  assign new_n4840_ = lo0442 & new_n4690_;
  assign new_n4841_ = lo0321 & new_n4693_;
  assign new_n4842_ = ~new_n4840_ & ~new_n4841_;
  assign new_n4843_ = lo0328 & new_n4681_;
  assign new_n4844_ = lo0459 & new_n4684_;
  assign new_n4845_ = ~new_n4843_ & ~new_n4844_;
  assign new_n4846_ = new_n4842_ & new_n4845_;
  assign new_n4847_ = lo0423 & new_n4684_;
  assign new_n4848_ = lo0348 & new_n4693_;
  assign new_n4849_ = ~new_n4847_ & ~new_n4848_;
  assign new_n4850_ = lo0398 & new_n4681_;
  assign new_n4851_ = lo0373 & new_n4690_;
  assign new_n4852_ = ~new_n4850_ & ~new_n4851_;
  assign new_n4853_ = new_n4849_ & new_n4852_;
  assign new_n4854_ = new_n4846_ & ~new_n4853_;
  assign new_n4855_ = ~new_n4846_ & new_n4853_;
  assign new_n4856_ = ~new_n4854_ & ~new_n4855_;
  assign new_n4857_ = new_n4839_ & ~new_n4856_;
  assign new_n4858_ = ~new_n4839_ & new_n4856_;
  assign new_n4859_ = ~new_n4857_ & ~new_n4858_;
  assign new_n4860_ = new_n4822_ & ~new_n4859_;
  assign new_n4861_ = ~new_n4822_ & new_n4859_;
  assign new_n4862_ = ~new_n4860_ & ~new_n4861_;
  assign new_n4863_ = new_n4785_ & ~new_n4862_;
  assign new_n4864_ = ~new_n4785_ & new_n4862_;
  assign new_n4865_ = ~new_n4863_ & ~new_n4864_;
  assign new_n4866_ = pi109 & ~new_n4865_;
  assign new_n4867_ = lo0433 & new_n4684_;
  assign new_n4868_ = lo0385 & new_n4690_;
  assign new_n4869_ = ~new_n4867_ & ~new_n4868_;
  assign new_n4870_ = lo0409 & new_n4681_;
  assign new_n4871_ = lo0360 & new_n4693_;
  assign new_n4872_ = ~new_n4870_ & ~new_n4871_;
  assign new_n4873_ = new_n4869_ & new_n4872_;
  assign new_n4874_ = lo0377 & new_n4690_;
  assign new_n4875_ = lo0462 & new_n4693_;
  assign new_n4876_ = ~new_n4874_ & ~new_n4875_;
  assign new_n4877_ = lo0318 & new_n4681_;
  assign new_n4878_ = lo0448 & new_n4684_;
  assign new_n4879_ = ~new_n4877_ & ~new_n4878_;
  assign new_n4880_ = new_n4876_ & new_n4879_;
  assign new_n4881_ = lo0381 & new_n4690_;
  assign new_n4882_ = lo0356 & new_n4693_;
  assign new_n4883_ = ~new_n4881_ & ~new_n4882_;
  assign new_n4884_ = lo0405 & new_n4681_;
  assign new_n4885_ = lo0445 & new_n4684_;
  assign new_n4886_ = ~new_n4884_ & ~new_n4885_;
  assign new_n4887_ = new_n4883_ & new_n4886_;
  assign new_n4888_ = new_n4880_ & ~new_n4887_;
  assign new_n4889_ = ~new_n4880_ & new_n4887_;
  assign new_n4890_ = ~new_n4888_ & ~new_n4889_;
  assign new_n4891_ = lo0326 & new_n4681_;
  assign new_n4892_ = lo0449 & new_n4684_;
  assign new_n4893_ = ~new_n4891_ & ~new_n4892_;
  assign new_n4894_ = lo0461 & new_n4693_;
  assign new_n4895_ = lo0439 & new_n4690_;
  assign new_n4896_ = ~new_n4894_ & ~new_n4895_;
  assign new_n4897_ = new_n4893_ & new_n4896_;
  assign new_n4898_ = lo0451 & new_n4684_;
  assign new_n4899_ = lo0353 & new_n4693_;
  assign new_n4900_ = ~new_n4898_ & ~new_n4899_;
  assign new_n4901_ = lo0325 & new_n4681_;
  assign new_n4902_ = lo0378 & new_n4690_;
  assign new_n4903_ = ~new_n4901_ & ~new_n4902_;
  assign new_n4904_ = new_n4900_ & new_n4903_;
  assign new_n4905_ = new_n4897_ & ~new_n4904_;
  assign new_n4906_ = ~new_n4897_ & new_n4904_;
  assign new_n4907_ = ~new_n4905_ & ~new_n4906_;
  assign new_n4908_ = new_n4890_ & ~new_n4907_;
  assign new_n4909_ = ~new_n4890_ & new_n4907_;
  assign new_n4910_ = ~new_n4908_ & ~new_n4909_;
  assign new_n4911_ = lo0382 & new_n4690_;
  assign new_n4912_ = lo0357 & new_n4693_;
  assign new_n4913_ = ~new_n4911_ & ~new_n4912_;
  assign new_n4914_ = lo0406 & new_n4681_;
  assign new_n4915_ = lo0430 & new_n4684_;
  assign new_n4916_ = ~new_n4914_ & ~new_n4915_;
  assign new_n4917_ = new_n4913_ & new_n4916_;
  assign new_n4918_ = lo0401 & new_n4681_;
  assign new_n4919_ = lo0351 & new_n4693_;
  assign new_n4920_ = ~new_n4918_ & ~new_n4919_;
  assign new_n4921_ = lo0426 & new_n4684_;
  assign new_n4922_ = lo0376 & new_n4690_;
  assign new_n4923_ = ~new_n4921_ & ~new_n4922_;
  assign new_n4924_ = new_n4920_ & new_n4923_;
  assign new_n4925_ = new_n4917_ & ~new_n4924_;
  assign new_n4926_ = ~new_n4917_ & new_n4924_;
  assign new_n4927_ = ~new_n4925_ & ~new_n4926_;
  assign new_n4928_ = lo0317 & new_n4690_;
  assign new_n4929_ = lo0352 & new_n4693_;
  assign new_n4930_ = ~new_n4928_ & ~new_n4929_;
  assign new_n4931_ = lo0402 & new_n4681_;
  assign new_n4932_ = lo0427 & new_n4684_;
  assign new_n4933_ = ~new_n4931_ & ~new_n4932_;
  assign new_n4934_ = new_n4930_ & new_n4933_;
  assign new_n4935_ = lo0379 & new_n4690_;
  assign new_n4936_ = lo0354 & new_n4693_;
  assign new_n4937_ = ~new_n4935_ & ~new_n4936_;
  assign new_n4938_ = lo0403 & new_n4681_;
  assign new_n4939_ = lo0428 & new_n4684_;
  assign new_n4940_ = ~new_n4938_ & ~new_n4939_;
  assign new_n4941_ = new_n4937_ & new_n4940_;
  assign new_n4942_ = new_n4934_ & ~new_n4941_;
  assign new_n4943_ = ~new_n4934_ & new_n4941_;
  assign new_n4944_ = ~new_n4942_ & ~new_n4943_;
  assign new_n4945_ = new_n4927_ & ~new_n4944_;
  assign new_n4946_ = ~new_n4927_ & new_n4944_;
  assign new_n4947_ = ~new_n4945_ & ~new_n4946_;
  assign new_n4948_ = new_n4910_ & ~new_n4947_;
  assign new_n4949_ = ~new_n4910_ & new_n4947_;
  assign new_n4950_ = ~new_n4948_ & ~new_n4949_;
  assign new_n4951_ = new_n4873_ & ~new_n4950_;
  assign new_n4952_ = ~new_n4873_ & new_n4950_;
  assign new_n4953_ = ~new_n4951_ & ~new_n4952_;
  assign new_n4954_ = pi110 & ~new_n4953_;
  assign new_n4955_ = lo0383 & new_n4690_;
  assign new_n4956_ = lo0358 & new_n4693_;
  assign new_n4957_ = ~new_n4955_ & ~new_n4956_;
  assign new_n4958_ = lo0407 & new_n4681_;
  assign new_n4959_ = lo0431 & new_n4684_;
  assign new_n4960_ = ~new_n4958_ & ~new_n4959_;
  assign new_n4961_ = new_n4957_ & new_n4960_;
  assign new_n4962_ = lo0364 & new_n4690_;
  assign new_n4963_ = lo0343 & new_n4693_;
  assign new_n4964_ = ~new_n4962_ & ~new_n4963_;
  assign new_n4965_ = lo0391 & new_n4681_;
  assign new_n4966_ = lo0415 & new_n4684_;
  assign new_n4967_ = ~new_n4965_ & ~new_n4966_;
  assign new_n4968_ = new_n4964_ & new_n4967_;
  assign new_n4969_ = lo0367 & new_n4690_;
  assign new_n4970_ = lo0345 & new_n4693_;
  assign new_n4971_ = ~new_n4969_ & ~new_n4970_;
  assign new_n4972_ = lo0392 & new_n4681_;
  assign new_n4973_ = lo0417 & new_n4684_;
  assign new_n4974_ = ~new_n4972_ & ~new_n4973_;
  assign new_n4975_ = new_n4971_ & new_n4974_;
  assign new_n4976_ = new_n4968_ & ~new_n4975_;
  assign new_n4977_ = ~new_n4968_ & new_n4975_;
  assign new_n4978_ = ~new_n4976_ & ~new_n4977_;
  assign new_n4979_ = lo0336 & new_n4690_;
  assign new_n4980_ = lo0362 & new_n4693_;
  assign new_n4981_ = ~new_n4979_ & ~new_n4980_;
  assign new_n4982_ = lo0463 & new_n4681_;
  assign new_n4983_ = lo0437 & new_n4684_;
  assign new_n4984_ = ~new_n4982_ & ~new_n4983_;
  assign new_n4985_ = new_n4981_ & new_n4984_;
  assign new_n4986_ = lo0447 & new_n4690_;
  assign new_n4987_ = lo0327 & new_n4693_;
  assign new_n4988_ = ~new_n4986_ & ~new_n4987_;
  assign new_n4989_ = lo0333 & new_n4681_;
  assign new_n4990_ = lo0453 & new_n4684_;
  assign new_n4991_ = ~new_n4989_ & ~new_n4990_;
  assign new_n4992_ = new_n4988_ & new_n4991_;
  assign new_n4993_ = new_n4985_ & ~new_n4992_;
  assign new_n4994_ = ~new_n4985_ & new_n4992_;
  assign new_n4995_ = ~new_n4993_ & ~new_n4994_;
  assign new_n4996_ = new_n4978_ & ~new_n4995_;
  assign new_n4997_ = ~new_n4978_ & new_n4995_;
  assign new_n4998_ = ~new_n4996_ & ~new_n4997_;
  assign new_n4999_ = lo0368 & new_n4690_;
  assign new_n5000_ = lo0346 & new_n4693_;
  assign new_n5001_ = ~new_n4999_ & ~new_n5000_;
  assign new_n5002_ = lo0393 & new_n4681_;
  assign new_n5003_ = lo0418 & new_n4684_;
  assign new_n5004_ = ~new_n5002_ & ~new_n5003_;
  assign new_n5005_ = new_n5001_ & new_n5004_;
  assign new_n5006_ = lo0389 & new_n4690_;
  assign new_n5007_ = lo0450 & new_n4693_;
  assign new_n5008_ = ~new_n5006_ & ~new_n5007_;
  assign new_n5009_ = lo0413 & new_n4681_;
  assign new_n5010_ = lo0438 & new_n4684_;
  assign new_n5011_ = ~new_n5009_ & ~new_n5010_;
  assign new_n5012_ = new_n5008_ & new_n5011_;
  assign new_n5013_ = new_n5005_ & ~new_n5012_;
  assign new_n5014_ = ~new_n5005_ & new_n5012_;
  assign new_n5015_ = ~new_n5013_ & ~new_n5014_;
  assign new_n5016_ = lo0365 & new_n4690_;
  assign new_n5017_ = lo0323 & new_n4693_;
  assign new_n5018_ = ~new_n5016_ & ~new_n5017_;
  assign new_n5019_ = lo0334 & new_n4681_;
  assign new_n5020_ = lo0464 & new_n4684_;
  assign new_n5021_ = ~new_n5019_ & ~new_n5020_;
  assign new_n5022_ = new_n5018_ & new_n5021_;
  assign new_n5023_ = lo0366 & new_n4690_;
  assign new_n5024_ = lo0344 & new_n4693_;
  assign new_n5025_ = ~new_n5023_ & ~new_n5024_;
  assign new_n5026_ = lo0335 & new_n4681_;
  assign new_n5027_ = lo0416 & new_n4684_;
  assign new_n5028_ = ~new_n5026_ & ~new_n5027_;
  assign new_n5029_ = new_n5025_ & new_n5028_;
  assign new_n5030_ = new_n5022_ & ~new_n5029_;
  assign new_n5031_ = ~new_n5022_ & new_n5029_;
  assign new_n5032_ = ~new_n5030_ & ~new_n5031_;
  assign new_n5033_ = new_n5015_ & ~new_n5032_;
  assign new_n5034_ = ~new_n5015_ & new_n5032_;
  assign new_n5035_ = ~new_n5033_ & ~new_n5034_;
  assign new_n5036_ = new_n4998_ & ~new_n5035_;
  assign new_n5037_ = ~new_n4998_ & new_n5035_;
  assign new_n5038_ = ~new_n5036_ & ~new_n5037_;
  assign new_n5039_ = new_n4961_ & ~new_n5038_;
  assign new_n5040_ = ~new_n4961_ & new_n5038_;
  assign new_n5041_ = ~new_n5039_ & ~new_n5040_;
  assign new_n5042_ = pi108 & ~new_n5041_;
  assign new_n5043_ = ~new_n4778_ & ~new_n4866_;
  assign new_n5044_ = ~new_n4954_ & new_n5043_;
  assign new_n5045_ = ~new_n5042_ & new_n5044_;
  assign new_n5046_ = new_n4678_ & ~new_n5045_;
  assign new_n5047_ = ~lo0098 & ~lo0567;
  assign new_n5048_ = new_n3673_ & ~new_n5047_;
  assign new_n5049_ = ~new_n5046_ & ~new_n5048_;
  assign new_n5050_ = ~pi072 & ~pi073;
  assign new_n5051_ = ~pi074 & new_n5050_;
  assign new_n5052_ = li0122 & new_n5049_;
  assign new_n5053_ = new_n5051_ & new_n5052_;
  assign new_n5054_ = pi072 & pi073;
  assign new_n5055_ = ~pi074 & new_n5054_;
  assign new_n5056_ = ~new_n5051_ & new_n5055_;
  assign new_n5057_ = ~lo0031 & new_n5056_;
  assign new_n5058_ = new_n3673_ & new_n5057_;
  assign li0031 = new_n5053_ | new_n5058_;
  assign new_n5060_ = ~new_n3979_ & ~new_n3985_;
  assign new_n5061_ = lo0032 & ~lo0314;
  assign new_n5062_ = ~lo0024 & lo0032;
  assign new_n5063_ = ~new_n5060_ & new_n5061_;
  assign new_n5064_ = new_n3940_ & new_n5062_;
  assign new_n5065_ = ~new_n5063_ & ~new_n5064_;
  assign new_n5066_ = lo0032 & ~lo0993;
  assign new_n5067_ = new_n3927_ & new_n5066_;
  assign new_n5068_ = new_n3953_ & new_n5062_;
  assign new_n5069_ = ~new_n5067_ & ~new_n5068_;
  assign new_n5070_ = new_n4424_ & new_n4653_;
  assign new_n5071_ = ~lo1076 & ~new_n4475_;
  assign new_n5072_ = lo0032 & new_n5071_;
  assign new_n5073_ = lo0032 & new_n4219_;
  assign new_n5074_ = lo0835 & ~li0583;
  assign new_n5075_ = ~new_n4427_ & ~new_n4428_;
  assign new_n5076_ = ~new_n4228_ & new_n5075_;
  assign new_n5077_ = lo0032 & li0583;
  assign new_n5078_ = new_n5073_ & ~new_n5074_;
  assign new_n5079_ = ~new_n5076_ & new_n5077_;
  assign new_n5080_ = ~new_n5078_ & ~new_n5079_;
  assign new_n5081_ = new_n4475_ & ~new_n5080_;
  assign new_n5082_ = lo1076 & ~new_n4475_;
  assign new_n5083_ = lo0786 & new_n5082_;
  assign new_n5084_ = lo0032 & new_n5083_;
  assign new_n5085_ = ~new_n5072_ & ~new_n5081_;
  assign new_n5086_ = ~new_n5084_ & new_n5085_;
  assign new_n5087_ = ~new_n4096_ & new_n5062_;
  assign new_n5088_ = lo0032 & ~new_n5062_;
  assign new_n5089_ = ~new_n5087_ & ~new_n5088_;
  assign new_n5090_ = new_n4023_ & ~new_n4091_;
  assign new_n5091_ = ~new_n5089_ & new_n5090_;
  assign new_n5092_ = new_n3746_ & new_n5061_;
  assign new_n5093_ = ~new_n5091_ & ~new_n5092_;
  assign new_n5094_ = new_n5070_ & ~new_n5086_;
  assign new_n5095_ = new_n5093_ & ~new_n5094_;
  assign new_n5096_ = ~new_n3589_ & ~new_n3735_;
  assign new_n5097_ = lo0032 & ~lo0841;
  assign new_n5098_ = new_n4020_ & new_n5062_;
  assign new_n5099_ = ~new_n5096_ & new_n5097_;
  assign new_n5100_ = ~new_n5098_ & ~new_n5099_;
  assign new_n5101_ = new_n5065_ & new_n5069_;
  assign new_n5102_ = new_n5095_ & new_n5101_;
  assign new_n5103_ = new_n5100_ & new_n5102_;
  assign new_n5104_ = ~new_n3862_ & ~new_n3867_;
  assign new_n5105_ = ~new_n3857_ & new_n5104_;
  assign new_n5106_ = new_n3804_ & new_n5062_;
  assign new_n5107_ = new_n3834_ & new_n5077_;
  assign new_n5108_ = new_n3678_ & new_n5107_;
  assign new_n5109_ = lo0479 & new_n3806_;
  assign new_n5110_ = new_n3809_ & new_n5109_;
  assign new_n5111_ = ~li0683 & new_n5110_;
  assign new_n5112_ = lo0841 & new_n5111_;
  assign new_n5113_ = lo0032 & new_n5112_;
  assign new_n5114_ = new_n3810_ & new_n5097_;
  assign new_n5115_ = ~new_n5106_ & ~new_n5108_;
  assign new_n5116_ = ~new_n5113_ & new_n5115_;
  assign new_n5117_ = ~new_n5114_ & new_n5116_;
  assign new_n5118_ = new_n5097_ & ~new_n5105_;
  assign new_n5119_ = new_n5117_ & ~new_n5118_;
  assign new_n5120_ = new_n3815_ & new_n5061_;
  assign new_n5121_ = new_n4088_ & new_n5062_;
  assign new_n5122_ = ~new_n5120_ & ~new_n5121_;
  assign new_n5123_ = ~lo1044 & new_n5061_;
  assign new_n5124_ = new_n3820_ & new_n5097_;
  assign new_n5125_ = new_n3870_ & new_n5123_;
  assign new_n5126_ = ~new_n5124_ & ~new_n5125_;
  assign new_n5127_ = ~new_n4069_ & new_n5062_;
  assign new_n5128_ = new_n5119_ & new_n5122_;
  assign new_n5129_ = new_n5126_ & new_n5128_;
  assign new_n5130_ = ~new_n5127_ & new_n5129_;
  assign new_n5131_ = ~lo0252 & new_n4647_;
  assign new_n5132_ = new_n3705_ & new_n4647_;
  assign new_n5133_ = ~new_n5131_ & new_n5132_;
  assign new_n5134_ = lo0252 & li0683;
  assign new_n5135_ = new_n5133_ & ~new_n5134_;
  assign new_n5136_ = lo0032 & new_n5135_;
  assign new_n5137_ = new_n3678_ & new_n4669_;
  assign new_n5138_ = new_n3890_ & ~new_n5137_;
  assign new_n5139_ = new_n3748_ & new_n5138_;
  assign new_n5140_ = new_n3678_ & new_n5139_;
  assign new_n5141_ = lo0032 & new_n5140_;
  assign new_n5142_ = new_n3786_ & new_n5062_;
  assign new_n5143_ = ~new_n5141_ & ~new_n5142_;
  assign new_n5144_ = new_n4041_ & new_n5062_;
  assign new_n5145_ = new_n5143_ & ~new_n5144_;
  assign new_n5146_ = lo0032 & lo1076;
  assign new_n5147_ = new_n3794_ & new_n5061_;
  assign new_n5148_ = new_n3763_ & new_n5097_;
  assign new_n5149_ = ~new_n5147_ & ~new_n5148_;
  assign new_n5150_ = new_n3914_ & new_n5061_;
  assign new_n5151_ = ~lo0137 & new_n4053_;
  assign new_n5152_ = lo0032 & ~new_n4632_;
  assign new_n5153_ = ~new_n5151_ & ~new_n5152_;
  assign new_n5154_ = new_n3777_ & ~new_n5153_;
  assign new_n5155_ = ~li0683 & ~new_n4669_;
  assign new_n5156_ = lo0032 & new_n5155_;
  assign new_n5157_ = new_n5154_ & ~new_n5155_;
  assign new_n5158_ = new_n3777_ & new_n5156_;
  assign new_n5159_ = ~new_n5157_ & ~new_n5158_;
  assign new_n5160_ = ~lo0024 & ~lo0032;
  assign new_n5161_ = new_n3780_ & ~new_n5160_;
  assign new_n5162_ = new_n3903_ & new_n5061_;
  assign new_n5163_ = ~new_n5161_ & ~new_n5162_;
  assign new_n5164_ = new_n5149_ & ~new_n5150_;
  assign new_n5165_ = new_n5159_ & new_n5164_;
  assign new_n5166_ = new_n5163_ & new_n5165_;
  assign new_n5167_ = new_n3773_ & new_n5146_;
  assign new_n5168_ = new_n5166_ & ~new_n5167_;
  assign new_n5169_ = lo0252 & ~new_n4647_;
  assign new_n5170_ = new_n4050_ & ~new_n5169_;
  assign new_n5171_ = new_n3655_ & new_n4647_;
  assign new_n5172_ = ~li0683 & ~new_n5171_;
  assign new_n5173_ = new_n5170_ & new_n5172_;
  assign new_n5174_ = ~lo0137 & new_n5173_;
  assign new_n5175_ = lo0024 & new_n5174_;
  assign new_n5176_ = new_n4050_ & new_n5062_;
  assign new_n5177_ = ~new_n5175_ & ~new_n5176_;
  assign new_n5178_ = ~new_n5136_ & new_n5145_;
  assign new_n5179_ = new_n5168_ & new_n5178_;
  assign new_n5180_ = new_n5177_ & new_n5179_;
  assign new_n5181_ = ~new_n3668_ & ~new_n3688_;
  assign new_n5182_ = ~lo0137 & ~new_n4647_;
  assign new_n5183_ = new_n5181_ & new_n5182_;
  assign new_n5184_ = ~lo0683 & new_n3678_;
  assign new_n5185_ = new_n4647_ & ~new_n5184_;
  assign new_n5186_ = ~new_n3688_ & new_n5185_;
  assign new_n5187_ = lo0032 & new_n5186_;
  assign new_n5188_ = ~new_n3668_ & new_n5187_;
  assign new_n5189_ = ~new_n5183_ & ~new_n5188_;
  assign new_n5190_ = ~new_n3689_ & ~new_n5189_;
  assign new_n5191_ = lo0032 & new_n3689_;
  assign new_n5192_ = ~new_n5190_ & ~new_n5191_;
  assign new_n5193_ = new_n3699_ & ~new_n5192_;
  assign new_n5194_ = lo0024 & new_n4135_;
  assign new_n5195_ = lo0032 & new_n5194_;
  assign new_n5196_ = ~new_n5062_ & ~new_n5195_;
  assign new_n5197_ = new_n3936_ & ~new_n5196_;
  assign new_n5198_ = new_n3625_ & new_n5062_;
  assign new_n5199_ = ~new_n5197_ & ~new_n5198_;
  assign new_n5200_ = ~new_n3725_ & ~new_n3931_;
  assign new_n5201_ = ~new_n3714_ & new_n5200_;
  assign new_n5202_ = new_n3969_ & new_n5097_;
  assign new_n5203_ = new_n5097_ & ~new_n5201_;
  assign new_n5204_ = ~new_n5202_ & ~new_n5203_;
  assign new_n5205_ = new_n4007_ & new_n5123_;
  assign new_n5206_ = new_n3948_ & new_n5062_;
  assign new_n5207_ = ~new_n5205_ & ~new_n5206_;
  assign new_n5208_ = new_n5199_ & new_n5204_;
  assign new_n5209_ = new_n5207_ & new_n5208_;
  assign new_n5210_ = lo0252 & li0583;
  assign new_n5211_ = lo0314 & ~new_n5210_;
  assign new_n5212_ = new_n4004_ & new_n5211_;
  assign new_n5213_ = lo0252 & ~lo0986;
  assign new_n5214_ = new_n4004_ & ~new_n5211_;
  assign new_n5215_ = new_n5212_ & new_n5213_;
  assign new_n5216_ = ~new_n5214_ & ~new_n5215_;
  assign new_n5217_ = lo0032 & ~new_n5216_;
  assign new_n5218_ = new_n4133_ & new_n5062_;
  assign new_n5219_ = ~new_n5217_ & ~new_n5218_;
  assign new_n5220_ = new_n3974_ & new_n5077_;
  assign new_n5221_ = ~new_n4135_ & new_n5220_;
  assign new_n5222_ = ~li0583 & ~new_n4053_;
  assign new_n5223_ = new_n3974_ & new_n5222_;
  assign new_n5224_ = lo0479 & new_n5223_;
  assign new_n5225_ = ~new_n4135_ & new_n5224_;
  assign new_n5226_ = lo0032 & new_n5225_;
  assign new_n5227_ = new_n5219_ & ~new_n5221_;
  assign new_n5228_ = ~new_n5226_ & new_n5227_;
  assign new_n5229_ = new_n5209_ & new_n5228_;
  assign new_n5230_ = new_n3678_ & new_n4647_;
  assign new_n5231_ = lo0032 & new_n4001_;
  assign new_n5232_ = new_n5230_ & new_n5231_;
  assign new_n5233_ = ~new_n5193_ & new_n5229_;
  assign new_n5234_ = ~new_n5232_ & new_n5233_;
  assign new_n5235_ = new_n5103_ & new_n5130_;
  assign new_n5236_ = new_n5180_ & new_n5235_;
  assign li0032 = ~new_n5234_ | ~new_n5236_;
  assign new_n5238_ = ~lo0979 & new_n4428_;
  assign new_n5239_ = ~new_n4421_ & new_n5238_;
  assign new_n5240_ = new_n4475_ & new_n5239_;
  assign new_n5241_ = new_n4135_ & new_n5240_;
  assign new_n5242_ = ~new_n4423_ & new_n5241_;
  assign new_n5243_ = new_n4653_ & new_n5242_;
  assign new_n5244_ = ~new_n3612_ & new_n4007_;
  assign new_n5245_ = ~new_n5243_ & ~new_n5244_;
  assign new_n5246_ = ~new_n4235_ & ~new_n5245_;
  assign new_n5247_ = ~new_n3612_ & new_n3870_;
  assign new_n5248_ = new_n4653_ & new_n5239_;
  assign new_n5249_ = ~new_n4423_ & new_n4528_;
  assign new_n5250_ = new_n4475_ & new_n5249_;
  assign new_n5251_ = new_n5248_ & new_n5250_;
  assign new_n5252_ = ~new_n5247_ & ~new_n5251_;
  assign new_n5253_ = new_n3633_ & new_n4543_;
  assign new_n5254_ = ~new_n3804_ & ~new_n3948_;
  assign new_n5255_ = ~new_n3786_ & new_n5254_;
  assign new_n5256_ = ~new_n3780_ & new_n5255_;
  assign new_n5257_ = ~new_n3953_ & new_n5256_;
  assign new_n5258_ = ~new_n4023_ & ~new_n5257_;
  assign new_n5259_ = ~new_n4535_ & ~new_n5258_;
  assign new_n5260_ = ~new_n4523_ & new_n5259_;
  assign new_n5261_ = new_n4347_ & new_n4543_;
  assign new_n5262_ = lo0164 & ~new_n3522_;
  assign new_n5263_ = lo0186 & new_n3522_;
  assign new_n5264_ = ~new_n5262_ & ~new_n5263_;
  assign new_n5265_ = new_n4543_ & new_n5264_;
  assign new_n5266_ = ~lo0038 & ~lo0059;
  assign new_n5267_ = ~lo0057 & new_n5266_;
  assign new_n5268_ = ~lo0054 & new_n5267_;
  assign new_n5269_ = ~lo0079 & ~lo0118;
  assign new_n5270_ = ~lo0033 & ~lo0139;
  assign new_n5271_ = ~lo0034 & new_n5270_;
  assign new_n5272_ = new_n5269_ & new_n5271_;
  assign new_n5273_ = ~lo0138 & new_n5272_;
  assign new_n5274_ = ~lo0195 & ~lo0196;
  assign li0841 = new_n5273_ & new_n5274_;
  assign new_n5276_ = ~lo0954 & ~li0841;
  assign new_n5277_ = ~lo0033 & ~new_n5276_;
  assign new_n5278_ = lo0033 & new_n5276_;
  assign new_n5279_ = ~new_n5277_ & ~new_n5278_;
  assign new_n5280_ = ~lo0040 & new_n3579_;
  assign new_n5281_ = ~new_n5279_ & new_n5280_;
  assign new_n5282_ = new_n5268_ & ~new_n5281_;
  assign new_n5283_ = ~new_n5265_ & ~new_n5268_;
  assign new_n5284_ = ~new_n5282_ & ~new_n5283_;
  assign new_n5285_ = ~lo0074 & ~new_n5284_;
  assign new_n5286_ = lo0074 & ~new_n5261_;
  assign new_n5287_ = ~new_n5285_ & ~new_n5286_;
  assign new_n5288_ = new_n5260_ & ~new_n5287_;
  assign new_n5289_ = new_n4523_ & new_n5259_;
  assign new_n5290_ = lo0183 & ~new_n3522_;
  assign new_n5291_ = lo0149 & ~lo0183;
  assign new_n5292_ = ~new_n5290_ & ~new_n5291_;
  assign new_n5293_ = new_n4543_ & new_n5292_;
  assign new_n5294_ = ~new_n5259_ & ~new_n5293_;
  assign new_n5295_ = ~new_n4557_ & new_n5289_;
  assign new_n5296_ = ~new_n5294_ & ~new_n5295_;
  assign new_n5297_ = ~lo0075 & ~lo0100;
  assign new_n5298_ = new_n5296_ & new_n5297_;
  assign new_n5299_ = lo0178 & ~new_n3522_;
  assign new_n5300_ = lo0157 & ~lo0178;
  assign new_n5301_ = ~new_n5299_ & ~new_n5300_;
  assign new_n5302_ = new_n4543_ & new_n5301_;
  assign new_n5303_ = ~new_n5293_ & ~new_n5302_;
  assign new_n5304_ = new_n5293_ & new_n5302_;
  assign new_n5305_ = ~new_n5303_ & ~new_n5304_;
  assign new_n5306_ = ~new_n5297_ & ~new_n5305_;
  assign new_n5307_ = new_n5252_ & ~new_n5306_;
  assign new_n5308_ = ~new_n5288_ & new_n5298_;
  assign new_n5309_ = new_n5307_ & ~new_n5308_;
  assign new_n5310_ = ~new_n5252_ & ~new_n5253_;
  assign new_n5311_ = ~new_n5309_ & ~new_n5310_;
  assign new_n5312_ = ~new_n3857_ & new_n3888_;
  assign new_n5313_ = ~new_n4637_ & ~new_n5312_;
  assign new_n5314_ = ~new_n4279_ & ~new_n5313_;
  assign new_n5315_ = ~new_n5311_ & new_n5313_;
  assign new_n5316_ = ~new_n5314_ & ~new_n5315_;
  assign new_n5317_ = ~new_n4543_ & ~new_n5313_;
  assign new_n5318_ = new_n5316_ & ~new_n5317_;
  assign new_n5319_ = new_n5245_ & ~new_n5318_;
  assign new_n5320_ = ~new_n5246_ & ~new_n5319_;
  assign new_n5321_ = ~new_n4543_ & ~new_n5245_;
  assign li0033 = ~new_n5320_ | new_n5321_;
  assign new_n5323_ = new_n3639_ & new_n4543_;
  assign new_n5324_ = new_n4330_ & new_n4543_;
  assign new_n5325_ = ~lo0033 & ~lo0034;
  assign new_n5326_ = lo0033 & lo0034;
  assign new_n5327_ = ~new_n5325_ & ~new_n5326_;
  assign new_n5328_ = new_n5276_ & ~new_n5327_;
  assign new_n5329_ = lo0034 & ~new_n5276_;
  assign new_n5330_ = ~new_n5328_ & ~new_n5329_;
  assign new_n5331_ = new_n5280_ & new_n5330_;
  assign new_n5332_ = new_n5268_ & ~new_n5331_;
  assign new_n5333_ = lo0167 & ~new_n3522_;
  assign new_n5334_ = lo0188 & new_n3522_;
  assign new_n5335_ = ~new_n5333_ & ~new_n5334_;
  assign new_n5336_ = new_n4543_ & new_n5335_;
  assign new_n5337_ = ~new_n5268_ & ~new_n5336_;
  assign new_n5338_ = ~new_n5332_ & ~new_n5337_;
  assign new_n5339_ = ~lo0074 & ~new_n5338_;
  assign new_n5340_ = lo0074 & ~new_n5324_;
  assign new_n5341_ = ~new_n5339_ & ~new_n5340_;
  assign new_n5342_ = new_n5260_ & ~new_n5341_;
  assign new_n5343_ = lo0140 & ~new_n3522_;
  assign new_n5344_ = ~lo0140 & lo0162;
  assign new_n5345_ = ~new_n5343_ & ~new_n5344_;
  assign new_n5346_ = new_n4543_ & new_n5345_;
  assign new_n5347_ = ~new_n5259_ & ~new_n5346_;
  assign new_n5348_ = ~new_n4548_ & new_n5289_;
  assign new_n5349_ = ~new_n5347_ & ~new_n5348_;
  assign new_n5350_ = new_n5297_ & new_n5349_;
  assign new_n5351_ = ~new_n5297_ & ~new_n5303_;
  assign new_n5352_ = ~new_n5297_ & new_n5303_;
  assign new_n5353_ = ~new_n4544_ & ~new_n5346_;
  assign new_n5354_ = new_n4544_ & new_n5346_;
  assign new_n5355_ = ~new_n5353_ & ~new_n5354_;
  assign new_n5356_ = new_n5351_ & new_n5355_;
  assign new_n5357_ = ~new_n5351_ & new_n5352_;
  assign new_n5358_ = ~new_n5356_ & ~new_n5357_;
  assign new_n5359_ = new_n5252_ & new_n5358_;
  assign new_n5360_ = ~new_n5342_ & new_n5350_;
  assign new_n5361_ = new_n5359_ & ~new_n5360_;
  assign new_n5362_ = ~new_n5252_ & ~new_n5323_;
  assign new_n5363_ = ~new_n5361_ & ~new_n5362_;
  assign new_n5364_ = new_n5313_ & ~new_n5363_;
  assign new_n5365_ = ~new_n3653_ & ~new_n5313_;
  assign new_n5366_ = ~new_n5244_ & ~new_n5365_;
  assign new_n5367_ = ~new_n5243_ & new_n5366_;
  assign new_n5368_ = ~new_n5317_ & new_n5367_;
  assign new_n5369_ = lo0177 & ~new_n3522_;
  assign new_n5370_ = lo0155 & ~lo0177;
  assign new_n5371_ = ~new_n5369_ & ~new_n5370_;
  assign new_n5372_ = ~new_n5245_ & new_n5371_;
  assign new_n5373_ = ~new_n5364_ & new_n5368_;
  assign new_n5374_ = ~new_n5372_ & ~new_n5373_;
  assign li0034 = new_n5321_ | new_n5374_;
  assign new_n5376_ = ~lo0024 & ~lo0035;
  assign new_n5377_ = lo0035 & ~lo0841;
  assign new_n5378_ = ~new_n3857_ & ~new_n3867_;
  assign new_n5379_ = new_n5377_ & ~new_n5378_;
  assign new_n5380_ = new_n4088_ & ~new_n5376_;
  assign new_n5381_ = ~new_n5379_ & ~new_n5380_;
  assign new_n5382_ = lo0035 & ~lo0314;
  assign new_n5383_ = new_n3618_ & ~new_n5376_;
  assign new_n5384_ = lo0035 & li0583;
  assign new_n5385_ = new_n3834_ & new_n5384_;
  assign new_n5386_ = new_n3678_ & new_n5385_;
  assign new_n5387_ = lo0035 & new_n5112_;
  assign new_n5388_ = new_n3810_ & new_n5377_;
  assign new_n5389_ = ~new_n5383_ & ~new_n5386_;
  assign new_n5390_ = ~new_n5387_ & new_n5389_;
  assign new_n5391_ = ~new_n5388_ & new_n5390_;
  assign new_n5392_ = new_n3815_ & new_n5382_;
  assign new_n5393_ = new_n5391_ & ~new_n5392_;
  assign new_n5394_ = ~new_n3804_ & ~new_n4068_;
  assign new_n5395_ = ~lo0024 & lo0035;
  assign new_n5396_ = ~new_n5394_ & new_n5395_;
  assign new_n5397_ = ~lo1044 & new_n5382_;
  assign new_n5398_ = new_n3820_ & new_n5377_;
  assign new_n5399_ = new_n3870_ & new_n5397_;
  assign new_n5400_ = ~new_n5398_ & ~new_n5399_;
  assign new_n5401_ = new_n5393_ & ~new_n5396_;
  assign new_n5402_ = new_n5400_ & new_n5401_;
  assign new_n5403_ = lo0035 & new_n3862_;
  assign new_n5404_ = new_n5402_ & ~new_n5403_;
  assign new_n5405_ = ~new_n4488_ & new_n5404_;
  assign new_n5406_ = lo0035 & new_n5071_;
  assign new_n5407_ = lo0035 & new_n4219_;
  assign new_n5408_ = ~new_n5074_ & new_n5407_;
  assign new_n5409_ = ~new_n5076_ & new_n5384_;
  assign new_n5410_ = ~new_n5408_ & ~new_n5409_;
  assign new_n5411_ = new_n4475_ & ~new_n5410_;
  assign new_n5412_ = lo0035 & new_n5083_;
  assign new_n5413_ = ~new_n5406_ & ~new_n5411_;
  assign new_n5414_ = ~new_n5412_ & new_n5413_;
  assign new_n5415_ = new_n3746_ & new_n5382_;
  assign new_n5416_ = ~new_n4096_ & ~new_n5376_;
  assign new_n5417_ = lo0035 & new_n5376_;
  assign new_n5418_ = ~new_n5416_ & ~new_n5417_;
  assign new_n5419_ = new_n5090_ & ~new_n5418_;
  assign new_n5420_ = ~new_n5415_ & ~new_n5419_;
  assign new_n5421_ = new_n5070_ & ~new_n5414_;
  assign new_n5422_ = new_n5420_ & ~new_n5421_;
  assign new_n5423_ = new_n4020_ & new_n5395_;
  assign new_n5424_ = ~new_n5096_ & new_n5377_;
  assign new_n5425_ = ~new_n5423_ & ~new_n5424_;
  assign new_n5426_ = new_n5381_ & new_n5405_;
  assign new_n5427_ = new_n5422_ & new_n5426_;
  assign new_n5428_ = new_n5425_ & new_n5427_;
  assign new_n5429_ = lo0137 & new_n5172_;
  assign new_n5430_ = ~new_n5169_ & ~new_n5429_;
  assign new_n5431_ = lo0024 & new_n4050_;
  assign new_n5432_ = ~new_n5430_ & new_n5431_;
  assign new_n5433_ = lo0035 & new_n5140_;
  assign new_n5434_ = new_n3786_ & new_n5395_;
  assign new_n5435_ = ~new_n5433_ & ~new_n5434_;
  assign new_n5436_ = ~new_n3888_ & new_n5435_;
  assign new_n5437_ = ~lo0035 & lo1076;
  assign new_n5438_ = new_n4050_ & new_n5395_;
  assign new_n5439_ = new_n4041_ & new_n5395_;
  assign new_n5440_ = ~new_n5438_ & ~new_n5439_;
  assign new_n5441_ = lo0035 & ~lo0993;
  assign new_n5442_ = new_n3927_ & new_n5441_;
  assign new_n5443_ = new_n3953_ & new_n5395_;
  assign new_n5444_ = ~new_n5442_ & ~new_n5443_;
  assign new_n5445_ = new_n5440_ & new_n5444_;
  assign new_n5446_ = new_n3773_ & ~new_n5437_;
  assign new_n5447_ = new_n5445_ & ~new_n5446_;
  assign new_n5448_ = ~new_n5432_ & new_n5436_;
  assign new_n5449_ = new_n5447_ & new_n5448_;
  assign new_n5450_ = lo0035 & ~new_n5216_;
  assign new_n5451_ = new_n4133_ & ~new_n5376_;
  assign new_n5452_ = ~new_n5450_ & ~new_n5451_;
  assign new_n5453_ = new_n3974_ & new_n5384_;
  assign new_n5454_ = ~new_n4135_ & new_n5453_;
  assign new_n5455_ = lo0035 & new_n5225_;
  assign new_n5456_ = new_n5452_ & ~new_n5454_;
  assign new_n5457_ = ~new_n5455_ & new_n5456_;
  assign new_n5458_ = new_n3948_ & new_n5395_;
  assign new_n5459_ = new_n5457_ & ~new_n5458_;
  assign new_n5460_ = ~new_n3903_ & ~new_n3914_;
  assign new_n5461_ = ~new_n5151_ & ~new_n5155_;
  assign new_n5462_ = ~lo0035 & ~new_n4632_;
  assign new_n5463_ = lo0035 & new_n5155_;
  assign new_n5464_ = new_n3777_ & new_n5463_;
  assign new_n5465_ = new_n3777_ & ~new_n5462_;
  assign new_n5466_ = new_n5461_ & new_n5465_;
  assign new_n5467_ = ~new_n5464_ & ~new_n5466_;
  assign new_n5468_ = new_n5382_ & ~new_n5460_;
  assign new_n5469_ = new_n5467_ & ~new_n5468_;
  assign new_n5470_ = new_n4007_ & new_n5397_;
  assign new_n5471_ = new_n3969_ & new_n5377_;
  assign new_n5472_ = ~new_n5470_ & ~new_n5471_;
  assign new_n5473_ = new_n3763_ & new_n5377_;
  assign new_n5474_ = new_n3780_ & new_n5395_;
  assign new_n5475_ = ~new_n5473_ & ~new_n5474_;
  assign new_n5476_ = new_n3794_ & new_n5382_;
  assign new_n5477_ = new_n5475_ & ~new_n5476_;
  assign new_n5478_ = new_n5459_ & new_n5469_;
  assign new_n5479_ = new_n5472_ & new_n5478_;
  assign new_n5480_ = new_n5477_ & new_n5479_;
  assign new_n5481_ = new_n5449_ & new_n5480_;
  assign new_n5482_ = new_n3940_ & new_n5395_;
  assign new_n5483_ = lo0035 & new_n5135_;
  assign new_n5484_ = ~new_n5482_ & ~new_n5483_;
  assign new_n5485_ = ~new_n5060_ & new_n5382_;
  assign new_n5486_ = new_n5484_ & ~new_n5485_;
  assign new_n5487_ = lo0035 & new_n5194_;
  assign new_n5488_ = ~new_n5395_ & ~new_n5487_;
  assign new_n5489_ = new_n3936_ & ~new_n5488_;
  assign new_n5490_ = new_n3625_ & new_n5395_;
  assign new_n5491_ = ~new_n5489_ & ~new_n5490_;
  assign new_n5492_ = ~new_n3668_ & ~new_n5182_;
  assign new_n5493_ = ~lo0035 & ~new_n5184_;
  assign new_n5494_ = new_n4647_ & new_n5493_;
  assign new_n5495_ = ~new_n3689_ & ~new_n5494_;
  assign new_n5496_ = new_n3688_ & ~new_n3689_;
  assign new_n5497_ = new_n5492_ & new_n5495_;
  assign new_n5498_ = ~new_n5496_ & ~new_n5497_;
  assign new_n5499_ = lo0035 & new_n3689_;
  assign new_n5500_ = new_n5498_ & ~new_n5499_;
  assign new_n5501_ = new_n3699_ & ~new_n5500_;
  assign new_n5502_ = new_n5491_ & ~new_n5501_;
  assign new_n5503_ = ~new_n5201_ & new_n5377_;
  assign new_n5504_ = new_n5502_ & ~new_n5503_;
  assign new_n5505_ = new_n4001_ & new_n5230_;
  assign new_n5506_ = lo0035 & new_n5505_;
  assign new_n5507_ = new_n5481_ & new_n5486_;
  assign new_n5508_ = new_n5504_ & new_n5507_;
  assign new_n5509_ = ~new_n5506_ & new_n5508_;
  assign li0035 = ~new_n5428_ | ~new_n5509_;
  assign new_n5511_ = lo0036 & ~lo0841;
  assign new_n5512_ = lo0036 & ~lo0314;
  assign new_n5513_ = new_n3746_ & new_n5512_;
  assign new_n5514_ = ~lo0024 & lo0036;
  assign new_n5515_ = new_n4020_ & new_n5514_;
  assign new_n5516_ = ~new_n5513_ & ~new_n5515_;
  assign new_n5517_ = ~new_n5096_ & new_n5511_;
  assign new_n5518_ = new_n5516_ & ~new_n5517_;
  assign new_n5519_ = new_n3804_ & new_n5514_;
  assign new_n5520_ = lo0036 & li0583;
  assign new_n5521_ = new_n3834_ & new_n5520_;
  assign new_n5522_ = new_n3678_ & new_n5521_;
  assign new_n5523_ = lo0036 & new_n5112_;
  assign new_n5524_ = new_n3810_ & new_n5511_;
  assign new_n5525_ = ~new_n5519_ & ~new_n5522_;
  assign new_n5526_ = ~new_n5523_ & new_n5525_;
  assign new_n5527_ = ~new_n5524_ & new_n5526_;
  assign new_n5528_ = ~new_n5105_ & new_n5511_;
  assign new_n5529_ = new_n5527_ & ~new_n5528_;
  assign new_n5530_ = new_n3815_ & new_n5512_;
  assign new_n5531_ = new_n4088_ & new_n5514_;
  assign new_n5532_ = ~new_n5530_ & ~new_n5531_;
  assign new_n5533_ = ~lo1044 & new_n5512_;
  assign new_n5534_ = new_n3820_ & new_n5511_;
  assign new_n5535_ = new_n3870_ & new_n5533_;
  assign new_n5536_ = ~new_n5534_ & ~new_n5535_;
  assign new_n5537_ = ~new_n4069_ & new_n5514_;
  assign new_n5538_ = new_n5536_ & ~new_n5537_;
  assign new_n5539_ = new_n5518_ & new_n5529_;
  assign new_n5540_ = new_n5532_ & new_n5539_;
  assign new_n5541_ = new_n5538_ & new_n5540_;
  assign new_n5542_ = lo0036 & new_n5071_;
  assign new_n5543_ = lo0036 & lo0786;
  assign new_n5544_ = ~new_n5076_ & new_n5520_;
  assign new_n5545_ = new_n4219_ & ~new_n5074_;
  assign new_n5546_ = lo0036 & new_n5545_;
  assign new_n5547_ = ~new_n5544_ & ~new_n5546_;
  assign new_n5548_ = new_n4475_ & ~new_n5547_;
  assign new_n5549_ = new_n5082_ & new_n5543_;
  assign new_n5550_ = ~new_n5548_ & ~new_n5549_;
  assign new_n5551_ = ~new_n5542_ & new_n5550_;
  assign new_n5552_ = new_n5070_ & ~new_n5551_;
  assign new_n5553_ = li0583 & new_n3753_;
  assign new_n5554_ = ~new_n4096_ & new_n5514_;
  assign new_n5555_ = lo0036 & ~new_n5514_;
  assign new_n5556_ = ~new_n5554_ & ~new_n5555_;
  assign new_n5557_ = new_n5090_ & ~new_n5556_;
  assign new_n5558_ = ~new_n5553_ & ~new_n5557_;
  assign new_n5559_ = ~new_n5552_ & new_n5558_;
  assign new_n5560_ = new_n5541_ & new_n5559_;
  assign new_n5561_ = new_n4050_ & new_n5514_;
  assign new_n5562_ = lo1076 & new_n3773_;
  assign new_n5563_ = lo0036 & new_n5562_;
  assign new_n5564_ = new_n3777_ & ~new_n5151_;
  assign new_n5565_ = ~new_n5155_ & new_n5564_;
  assign new_n5566_ = lo0036 & new_n5155_;
  assign new_n5567_ = new_n3777_ & new_n5566_;
  assign new_n5568_ = lo0036 & ~new_n4632_;
  assign new_n5569_ = new_n5565_ & new_n5568_;
  assign new_n5570_ = ~new_n5567_ & ~new_n5569_;
  assign new_n5571_ = ~new_n5460_ & new_n5512_;
  assign new_n5572_ = new_n5570_ & ~new_n5571_;
  assign new_n5573_ = new_n3763_ & new_n5511_;
  assign new_n5574_ = new_n3780_ & new_n5514_;
  assign new_n5575_ = ~new_n5573_ & ~new_n5574_;
  assign new_n5576_ = new_n3794_ & new_n5512_;
  assign new_n5577_ = new_n5575_ & ~new_n5576_;
  assign new_n5578_ = ~new_n5561_ & ~new_n5563_;
  assign new_n5579_ = new_n5572_ & new_n5578_;
  assign new_n5580_ = new_n5577_ & new_n5579_;
  assign new_n5581_ = new_n4041_ & new_n5514_;
  assign new_n5582_ = new_n5580_ & ~new_n5581_;
  assign new_n5583_ = lo0036 & new_n3678_;
  assign new_n5584_ = new_n3786_ & new_n5514_;
  assign new_n5585_ = new_n5139_ & new_n5583_;
  assign new_n5586_ = ~new_n5584_ & ~new_n5585_;
  assign new_n5587_ = new_n4007_ & new_n5533_;
  assign new_n5588_ = new_n3969_ & new_n5511_;
  assign new_n5589_ = ~new_n5587_ & ~new_n5588_;
  assign new_n5590_ = lo0036 & ~new_n5216_;
  assign new_n5591_ = new_n4133_ & new_n5514_;
  assign new_n5592_ = ~new_n5590_ & ~new_n5591_;
  assign new_n5593_ = new_n3974_ & new_n5520_;
  assign new_n5594_ = ~new_n4135_ & new_n5593_;
  assign new_n5595_ = lo0036 & new_n5225_;
  assign new_n5596_ = new_n5592_ & ~new_n5594_;
  assign new_n5597_ = ~new_n5595_ & new_n5596_;
  assign new_n5598_ = new_n3948_ & new_n5514_;
  assign new_n5599_ = new_n5597_ & ~new_n5598_;
  assign new_n5600_ = new_n5582_ & new_n5586_;
  assign new_n5601_ = new_n5589_ & new_n5600_;
  assign new_n5602_ = new_n5599_ & new_n5601_;
  assign new_n5603_ = lo0036 & new_n5505_;
  assign new_n5604_ = lo0036 & new_n5135_;
  assign new_n5605_ = ~new_n3688_ & new_n3699_;
  assign new_n5606_ = ~new_n3689_ & new_n5605_;
  assign new_n5607_ = ~new_n3668_ & new_n5606_;
  assign new_n5608_ = new_n4647_ & new_n5607_;
  assign new_n5609_ = lo0036 & new_n5608_;
  assign new_n5610_ = ~new_n5184_ & new_n5609_;
  assign new_n5611_ = lo0036 & li0683;
  assign new_n5612_ = ~li0583 & ~new_n5611_;
  assign new_n5613_ = new_n4631_ & ~new_n5612_;
  assign new_n5614_ = new_n3936_ & new_n5514_;
  assign new_n5615_ = ~new_n5613_ & ~new_n5614_;
  assign new_n5616_ = new_n3625_ & new_n5514_;
  assign new_n5617_ = lo0036 & new_n3706_;
  assign new_n5618_ = ~new_n5610_ & new_n5615_;
  assign new_n5619_ = ~new_n5616_ & new_n5618_;
  assign new_n5620_ = ~new_n5617_ & new_n5619_;
  assign new_n5621_ = ~new_n5201_ & new_n5511_;
  assign new_n5622_ = new_n5620_ & ~new_n5621_;
  assign new_n5623_ = ~new_n5603_ & ~new_n5604_;
  assign new_n5624_ = new_n5622_ & new_n5623_;
  assign new_n5625_ = new_n5602_ & new_n5624_;
  assign new_n5626_ = ~new_n5060_ & new_n5512_;
  assign new_n5627_ = new_n3940_ & new_n5514_;
  assign new_n5628_ = ~new_n5626_ & ~new_n5627_;
  assign new_n5629_ = lo0036 & ~lo0993;
  assign new_n5630_ = new_n3927_ & new_n5629_;
  assign new_n5631_ = new_n3953_ & new_n5514_;
  assign new_n5632_ = ~new_n5630_ & ~new_n5631_;
  assign new_n5633_ = new_n5628_ & new_n5632_;
  assign new_n5634_ = new_n5560_ & new_n5625_;
  assign li0036 = ~new_n5633_ | ~new_n5634_;
  assign new_n5636_ = ~lo0024 & lo0038;
  assign new_n5637_ = new_n4050_ & new_n5636_;
  assign new_n5638_ = lo0038 & new_n5562_;
  assign new_n5639_ = lo0038 & ~lo0314;
  assign new_n5640_ = lo0038 & new_n5155_;
  assign new_n5641_ = new_n3777_ & new_n5640_;
  assign new_n5642_ = lo0038 & ~new_n4632_;
  assign new_n5643_ = new_n5565_ & new_n5642_;
  assign new_n5644_ = ~new_n5641_ & ~new_n5643_;
  assign new_n5645_ = ~new_n5460_ & new_n5639_;
  assign new_n5646_ = new_n5644_ & ~new_n5645_;
  assign new_n5647_ = lo0038 & ~lo0841;
  assign new_n5648_ = new_n3763_ & new_n5647_;
  assign new_n5649_ = new_n3780_ & new_n5636_;
  assign new_n5650_ = ~new_n5648_ & ~new_n5649_;
  assign new_n5651_ = new_n3794_ & new_n5639_;
  assign new_n5652_ = new_n5650_ & ~new_n5651_;
  assign new_n5653_ = ~new_n5637_ & ~new_n5638_;
  assign new_n5654_ = new_n5646_ & new_n5653_;
  assign new_n5655_ = new_n5652_ & new_n5654_;
  assign new_n5656_ = new_n4041_ & new_n5636_;
  assign new_n5657_ = new_n5655_ & ~new_n5656_;
  assign new_n5658_ = lo0038 & new_n3706_;
  assign new_n5659_ = lo0038 & new_n5194_;
  assign new_n5660_ = ~new_n5636_ & ~new_n5659_;
  assign new_n5661_ = new_n3936_ & ~new_n5660_;
  assign new_n5662_ = ~lo0038 & ~lo0841;
  assign new_n5663_ = new_n3714_ & ~new_n5662_;
  assign new_n5664_ = new_n3725_ & new_n5647_;
  assign new_n5665_ = ~new_n5663_ & ~new_n5664_;
  assign new_n5666_ = ~new_n5658_ & ~new_n5661_;
  assign new_n5667_ = new_n5665_ & new_n5666_;
  assign new_n5668_ = ~new_n5060_ & new_n5639_;
  assign new_n5669_ = new_n3940_ & new_n5636_;
  assign new_n5670_ = ~new_n5668_ & ~new_n5669_;
  assign new_n5671_ = ~lo0993 & new_n3927_;
  assign new_n5672_ = lo0038 & new_n5671_;
  assign new_n5673_ = new_n3953_ & new_n5636_;
  assign new_n5674_ = new_n5670_ & ~new_n5672_;
  assign new_n5675_ = ~new_n5673_ & new_n5674_;
  assign new_n5676_ = new_n5667_ & new_n5675_;
  assign new_n5677_ = new_n5657_ & new_n5676_;
  assign new_n5678_ = lo0038 & new_n5230_;
  assign new_n5679_ = lo0038 & new_n3678_;
  assign new_n5680_ = new_n3786_ & new_n5636_;
  assign new_n5681_ = new_n5139_ & new_n5679_;
  assign new_n5682_ = ~new_n5680_ & ~new_n5681_;
  assign new_n5683_ = lo0038 & ~new_n5134_;
  assign new_n5684_ = new_n5133_ & new_n5683_;
  assign new_n5685_ = ~lo1044 & new_n5639_;
  assign new_n5686_ = new_n4007_ & new_n5685_;
  assign new_n5687_ = new_n3948_ & new_n5636_;
  assign new_n5688_ = ~new_n5686_ & ~new_n5687_;
  assign new_n5689_ = new_n3931_ & new_n5647_;
  assign new_n5690_ = new_n3625_ & new_n5636_;
  assign new_n5691_ = ~new_n5689_ & ~new_n5690_;
  assign new_n5692_ = new_n5682_ & ~new_n5684_;
  assign new_n5693_ = new_n5688_ & new_n5692_;
  assign new_n5694_ = new_n5691_ & new_n5693_;
  assign new_n5695_ = new_n4001_ & new_n5678_;
  assign new_n5696_ = new_n5694_ & ~new_n5695_;
  assign new_n5697_ = lo0038 & ~new_n5216_;
  assign new_n5698_ = new_n3969_ & new_n5647_;
  assign new_n5699_ = ~new_n5697_ & ~new_n5698_;
  assign new_n5700_ = lo0038 & li0583;
  assign new_n5701_ = new_n3974_ & new_n5700_;
  assign new_n5702_ = ~new_n4135_ & new_n5701_;
  assign new_n5703_ = lo0038 & new_n5225_;
  assign new_n5704_ = new_n5699_ & ~new_n5702_;
  assign new_n5705_ = ~new_n5703_ & new_n5704_;
  assign new_n5706_ = new_n4133_ & new_n5636_;
  assign new_n5707_ = new_n5705_ & ~new_n5706_;
  assign new_n5708_ = ~new_n5184_ & new_n5608_;
  assign new_n5709_ = lo0038 & new_n5708_;
  assign new_n5710_ = new_n5696_ & new_n5707_;
  assign new_n5711_ = ~new_n5709_ & new_n5710_;
  assign new_n5712_ = new_n5677_ & new_n5711_;
  assign new_n5713_ = lo0332 & lo0841;
  assign new_n5714_ = ~new_n5647_ & ~new_n5713_;
  assign new_n5715_ = lo0038 & new_n5071_;
  assign new_n5716_ = lo0038 & lo0786;
  assign new_n5717_ = ~new_n5076_ & new_n5700_;
  assign new_n5718_ = lo0038 & new_n5545_;
  assign new_n5719_ = ~new_n5717_ & ~new_n5718_;
  assign new_n5720_ = new_n4475_ & ~new_n5719_;
  assign new_n5721_ = new_n5082_ & new_n5716_;
  assign new_n5722_ = ~new_n5720_ & ~new_n5721_;
  assign new_n5723_ = ~new_n5715_ & new_n5722_;
  assign new_n5724_ = new_n4653_ & ~new_n5723_;
  assign new_n5725_ = ~new_n4096_ & new_n5636_;
  assign new_n5726_ = lo0038 & ~new_n5636_;
  assign new_n5727_ = ~new_n5725_ & ~new_n5726_;
  assign new_n5728_ = new_n4424_ & new_n5724_;
  assign new_n5729_ = new_n5090_ & ~new_n5727_;
  assign new_n5730_ = ~new_n5728_ & ~new_n5729_;
  assign new_n5731_ = new_n3589_ & ~new_n5714_;
  assign new_n5732_ = new_n5730_ & ~new_n5731_;
  assign new_n5733_ = new_n3746_ & new_n5639_;
  assign new_n5734_ = new_n5732_ & ~new_n5733_;
  assign new_n5735_ = new_n4020_ & new_n5636_;
  assign new_n5736_ = new_n3735_ & new_n5647_;
  assign new_n5737_ = ~new_n5735_ & ~new_n5736_;
  assign new_n5738_ = new_n3862_ & new_n5647_;
  assign new_n5739_ = new_n4088_ & new_n5636_;
  assign new_n5740_ = ~new_n5738_ & ~new_n5739_;
  assign new_n5741_ = new_n3867_ & new_n5647_;
  assign new_n5742_ = new_n3815_ & new_n5639_;
  assign new_n5743_ = ~new_n5741_ & ~new_n5742_;
  assign new_n5744_ = new_n3618_ & new_n5636_;
  assign new_n5745_ = new_n3870_ & new_n5685_;
  assign new_n5746_ = ~new_n5744_ & ~new_n5745_;
  assign new_n5747_ = ~new_n5394_ & new_n5636_;
  assign new_n5748_ = new_n5746_ & ~new_n5747_;
  assign new_n5749_ = lo0038 & lo0841;
  assign new_n5750_ = new_n3810_ & new_n5647_;
  assign new_n5751_ = new_n5111_ & new_n5749_;
  assign new_n5752_ = ~new_n5750_ & ~new_n5751_;
  assign new_n5753_ = new_n3678_ & new_n5700_;
  assign new_n5754_ = new_n3834_ & new_n5753_;
  assign new_n5755_ = new_n3820_ & new_n5647_;
  assign new_n5756_ = ~new_n5754_ & ~new_n5755_;
  assign new_n5757_ = new_n5743_ & new_n5748_;
  assign new_n5758_ = new_n5752_ & new_n5757_;
  assign new_n5759_ = new_n5756_ & new_n5758_;
  assign new_n5760_ = new_n3857_ & new_n5647_;
  assign new_n5761_ = new_n5759_ & ~new_n5760_;
  assign new_n5762_ = new_n5734_ & new_n5737_;
  assign new_n5763_ = new_n5740_ & new_n5762_;
  assign new_n5764_ = new_n5761_ & new_n5763_;
  assign li0038 = ~new_n5712_ | ~new_n5764_;
  assign new_n5766_ = lo0039 & ~lo0841;
  assign new_n5767_ = ~lo0024 & lo0039;
  assign new_n5768_ = new_n4020_ & new_n5767_;
  assign new_n5769_ = ~new_n5096_ & new_n5766_;
  assign new_n5770_ = ~new_n5768_ & ~new_n5769_;
  assign new_n5771_ = lo0039 & new_n5071_;
  assign new_n5772_ = lo0039 & lo0786;
  assign new_n5773_ = lo0039 & li0583;
  assign new_n5774_ = ~new_n5076_ & new_n5773_;
  assign new_n5775_ = lo0039 & new_n5545_;
  assign new_n5776_ = ~new_n5774_ & ~new_n5775_;
  assign new_n5777_ = new_n4475_ & ~new_n5776_;
  assign new_n5778_ = new_n5082_ & new_n5772_;
  assign new_n5779_ = ~new_n5777_ & ~new_n5778_;
  assign new_n5780_ = ~new_n5771_ & new_n5779_;
  assign new_n5781_ = new_n4653_ & ~new_n5780_;
  assign new_n5782_ = lo0039 & ~lo0314;
  assign new_n5783_ = new_n4424_ & new_n5781_;
  assign new_n5784_ = new_n3746_ & new_n5782_;
  assign new_n5785_ = ~new_n5783_ & ~new_n5784_;
  assign new_n5786_ = ~new_n4096_ & new_n5767_;
  assign new_n5787_ = lo0039 & ~new_n5767_;
  assign new_n5788_ = ~new_n5786_ & ~new_n5787_;
  assign new_n5789_ = new_n4023_ & ~new_n5788_;
  assign new_n5790_ = new_n5770_ & new_n5785_;
  assign new_n5791_ = ~new_n4498_ & new_n5790_;
  assign new_n5792_ = ~new_n5789_ & new_n5791_;
  assign new_n5793_ = lo0039 & ~lo0993;
  assign new_n5794_ = new_n3927_ & new_n5793_;
  assign new_n5795_ = new_n3953_ & new_n5767_;
  assign new_n5796_ = ~new_n5794_ & ~new_n5795_;
  assign new_n5797_ = ~lo1044 & new_n5782_;
  assign new_n5798_ = new_n4007_ & new_n5797_;
  assign new_n5799_ = new_n3969_ & new_n5766_;
  assign new_n5800_ = ~new_n5798_ & ~new_n5799_;
  assign new_n5801_ = ~new_n3996_ & new_n5800_;
  assign new_n5802_ = new_n4133_ & new_n5767_;
  assign new_n5803_ = ~lo0039 & new_n5213_;
  assign new_n5804_ = new_n5212_ & ~new_n5803_;
  assign new_n5805_ = lo0039 & ~new_n5211_;
  assign new_n5806_ = new_n4004_ & new_n5805_;
  assign new_n5807_ = ~new_n5802_ & ~new_n5804_;
  assign new_n5808_ = ~new_n5806_ & new_n5807_;
  assign new_n5809_ = ~new_n4135_ & new_n5773_;
  assign new_n5810_ = new_n3974_ & new_n5809_;
  assign new_n5811_ = lo0039 & ~new_n4135_;
  assign new_n5812_ = new_n5224_ & new_n5811_;
  assign new_n5813_ = ~new_n5810_ & ~new_n5812_;
  assign new_n5814_ = new_n5808_ & new_n5813_;
  assign new_n5815_ = ~new_n3668_ & ~new_n3689_;
  assign new_n5816_ = ~new_n3688_ & new_n5815_;
  assign new_n5817_ = new_n3699_ & new_n5816_;
  assign new_n5818_ = new_n4647_ & new_n5817_;
  assign new_n5819_ = lo0039 & new_n5818_;
  assign new_n5820_ = ~new_n5184_ & new_n5819_;
  assign new_n5821_ = ~lo0039 & ~lo0841;
  assign new_n5822_ = lo0039 & new_n5194_;
  assign new_n5823_ = ~new_n5767_ & ~new_n5822_;
  assign new_n5824_ = new_n3936_ & ~new_n5823_;
  assign new_n5825_ = new_n3725_ & ~new_n5821_;
  assign new_n5826_ = ~new_n5824_ & ~new_n5825_;
  assign new_n5827_ = ~new_n3714_ & ~new_n3931_;
  assign new_n5828_ = new_n5766_ & ~new_n5827_;
  assign new_n5829_ = new_n3625_ & new_n5767_;
  assign new_n5830_ = ~new_n5828_ & ~new_n5829_;
  assign new_n5831_ = lo0039 & new_n3706_;
  assign new_n5832_ = ~new_n5820_ & new_n5826_;
  assign new_n5833_ = new_n5830_ & new_n5832_;
  assign new_n5834_ = ~new_n5831_ & new_n5833_;
  assign new_n5835_ = new_n3948_ & new_n5767_;
  assign new_n5836_ = new_n5834_ & ~new_n5835_;
  assign new_n5837_ = new_n5796_ & new_n5801_;
  assign new_n5838_ = new_n5814_ & new_n5837_;
  assign new_n5839_ = new_n5836_ & new_n5838_;
  assign new_n5840_ = new_n5792_ & new_n5839_;
  assign new_n5841_ = ~new_n3863_ & new_n5766_;
  assign new_n5842_ = new_n4088_ & new_n5767_;
  assign new_n5843_ = ~new_n5841_ & ~new_n5842_;
  assign new_n5844_ = new_n3867_ & ~new_n5821_;
  assign new_n5845_ = new_n3815_ & new_n5782_;
  assign new_n5846_ = ~new_n5844_ & ~new_n5845_;
  assign new_n5847_ = new_n3820_ & new_n5766_;
  assign new_n5848_ = new_n3870_ & new_n5797_;
  assign new_n5849_ = ~new_n5847_ & ~new_n5848_;
  assign new_n5850_ = ~new_n4069_ & new_n5767_;
  assign new_n5851_ = new_n5849_ & ~new_n5850_;
  assign new_n5852_ = new_n3834_ & new_n5773_;
  assign new_n5853_ = new_n3678_ & new_n5852_;
  assign new_n5854_ = new_n3804_ & new_n5767_;
  assign new_n5855_ = ~new_n5853_ & ~new_n5854_;
  assign new_n5856_ = lo0039 & new_n5112_;
  assign new_n5857_ = new_n3810_ & new_n5766_;
  assign new_n5858_ = ~new_n5856_ & ~new_n5857_;
  assign new_n5859_ = new_n5855_ & new_n5858_;
  assign new_n5860_ = new_n5843_ & new_n5846_;
  assign new_n5861_ = new_n5851_ & new_n5860_;
  assign new_n5862_ = new_n5859_ & new_n5861_;
  assign new_n5863_ = new_n3940_ & new_n5767_;
  assign new_n5864_ = lo0039 & new_n5135_;
  assign new_n5865_ = ~new_n5863_ & ~new_n5864_;
  assign new_n5866_ = ~new_n5060_ & new_n5782_;
  assign new_n5867_ = new_n5865_ & ~new_n5866_;
  assign new_n5868_ = lo0039 & new_n5505_;
  assign new_n5869_ = lo0039 & new_n3678_;
  assign new_n5870_ = new_n3786_ & new_n5767_;
  assign new_n5871_ = new_n5139_ & new_n5869_;
  assign new_n5872_ = ~new_n5870_ & ~new_n5871_;
  assign new_n5873_ = new_n3780_ & new_n5767_;
  assign new_n5874_ = lo0039 & new_n5155_;
  assign new_n5875_ = new_n3777_ & new_n5874_;
  assign new_n5876_ = lo0039 & ~new_n4632_;
  assign new_n5877_ = new_n5565_ & new_n5876_;
  assign new_n5878_ = ~new_n5875_ & ~new_n5877_;
  assign new_n5879_ = ~new_n5873_ & new_n5878_;
  assign new_n5880_ = new_n3763_ & new_n5766_;
  assign new_n5881_ = lo0039 & new_n3773_;
  assign new_n5882_ = lo1076 & new_n5881_;
  assign new_n5883_ = new_n3794_ & new_n5782_;
  assign new_n5884_ = ~new_n5460_ & new_n5782_;
  assign new_n5885_ = ~new_n5883_ & ~new_n5884_;
  assign new_n5886_ = ~new_n5882_ & new_n5885_;
  assign new_n5887_ = new_n4050_ & new_n5767_;
  assign new_n5888_ = new_n5886_ & ~new_n5887_;
  assign new_n5889_ = ~new_n5880_ & new_n5888_;
  assign new_n5890_ = new_n5879_ & new_n5889_;
  assign new_n5891_ = new_n4041_ & new_n5767_;
  assign new_n5892_ = new_n5890_ & ~new_n5891_;
  assign new_n5893_ = new_n5867_ & ~new_n5868_;
  assign new_n5894_ = new_n5872_ & new_n5893_;
  assign new_n5895_ = new_n5892_ & new_n5894_;
  assign new_n5896_ = new_n5862_ & new_n5895_;
  assign li0039 = ~new_n5840_ | ~new_n5896_;
  assign new_n5898_ = lo0040 & new_n3706_;
  assign new_n5899_ = lo0040 & new_n4135_;
  assign new_n5900_ = ~lo0024 & lo0040;
  assign new_n5901_ = lo0024 & new_n5899_;
  assign new_n5902_ = ~new_n5900_ & ~new_n5901_;
  assign new_n5903_ = new_n3936_ & ~new_n5902_;
  assign new_n5904_ = lo0040 & ~lo0841;
  assign new_n5905_ = new_n3725_ & new_n5904_;
  assign new_n5906_ = new_n3625_ & new_n5900_;
  assign new_n5907_ = ~new_n5905_ & ~new_n5906_;
  assign new_n5908_ = ~new_n5827_ & new_n5904_;
  assign new_n5909_ = new_n5907_ & ~new_n5908_;
  assign new_n5910_ = ~new_n5898_ & ~new_n5903_;
  assign new_n5911_ = new_n5909_ & new_n5910_;
  assign new_n5912_ = ~new_n4018_ & new_n5911_;
  assign new_n5913_ = lo0040 & ~lo0314;
  assign new_n5914_ = ~new_n5060_ & new_n5913_;
  assign new_n5915_ = new_n3940_ & new_n5900_;
  assign new_n5916_ = ~new_n5914_ & ~new_n5915_;
  assign new_n5917_ = new_n3953_ & new_n5900_;
  assign new_n5918_ = lo0040 & new_n5671_;
  assign new_n5919_ = new_n5916_ & ~new_n5917_;
  assign new_n5920_ = ~new_n5918_ & new_n5919_;
  assign new_n5921_ = new_n5912_ & new_n5920_;
  assign new_n5922_ = lo0040 & new_n3678_;
  assign new_n5923_ = new_n3786_ & new_n5900_;
  assign new_n5924_ = new_n5139_ & new_n5922_;
  assign new_n5925_ = ~new_n5923_ & ~new_n5924_;
  assign new_n5926_ = lo0040 & new_n5135_;
  assign new_n5927_ = ~lo1044 & new_n5913_;
  assign new_n5928_ = new_n4007_ & new_n5927_;
  assign new_n5929_ = new_n3969_ & new_n5904_;
  assign new_n5930_ = ~new_n5928_ & ~new_n5929_;
  assign new_n5931_ = new_n5921_ & new_n5925_;
  assign new_n5932_ = ~new_n5926_ & new_n5931_;
  assign new_n5933_ = new_n5930_ & new_n5932_;
  assign new_n5934_ = new_n4050_ & new_n5900_;
  assign new_n5935_ = lo0040 & new_n5562_;
  assign new_n5936_ = lo0040 & new_n5155_;
  assign new_n5937_ = new_n3777_ & new_n5936_;
  assign new_n5938_ = lo0040 & ~new_n4632_;
  assign new_n5939_ = new_n5565_ & new_n5938_;
  assign new_n5940_ = ~new_n5937_ & ~new_n5939_;
  assign new_n5941_ = ~new_n5460_ & new_n5913_;
  assign new_n5942_ = new_n5940_ & ~new_n5941_;
  assign new_n5943_ = new_n3763_ & new_n5904_;
  assign new_n5944_ = new_n3780_ & new_n5900_;
  assign new_n5945_ = ~new_n5943_ & ~new_n5944_;
  assign new_n5946_ = new_n3794_ & new_n5913_;
  assign new_n5947_ = new_n5945_ & ~new_n5946_;
  assign new_n5948_ = ~new_n5934_ & ~new_n5935_;
  assign new_n5949_ = new_n5942_ & new_n5948_;
  assign new_n5950_ = new_n5947_ & new_n5949_;
  assign new_n5951_ = new_n4041_ & new_n5900_;
  assign new_n5952_ = new_n5950_ & ~new_n5951_;
  assign new_n5953_ = lo0040 & ~new_n5216_;
  assign new_n5954_ = new_n4133_ & new_n5900_;
  assign new_n5955_ = ~new_n5953_ & ~new_n5954_;
  assign new_n5956_ = lo0040 & li0583;
  assign new_n5957_ = new_n3974_ & new_n5956_;
  assign new_n5958_ = ~new_n4135_ & new_n5957_;
  assign new_n5959_ = lo0040 & new_n5225_;
  assign new_n5960_ = new_n5955_ & ~new_n5958_;
  assign new_n5961_ = ~new_n5959_ & new_n5960_;
  assign new_n5962_ = new_n3948_ & new_n5900_;
  assign new_n5963_ = new_n5961_ & ~new_n5962_;
  assign new_n5964_ = lo0040 & new_n5708_;
  assign new_n5965_ = lo0040 & new_n5230_;
  assign new_n5966_ = new_n4001_ & new_n5965_;
  assign new_n5967_ = new_n5952_ & new_n5963_;
  assign new_n5968_ = ~new_n5964_ & new_n5967_;
  assign new_n5969_ = ~new_n5966_ & new_n5968_;
  assign new_n5970_ = new_n5933_ & new_n5969_;
  assign new_n5971_ = new_n4020_ & new_n5900_;
  assign new_n5972_ = ~new_n5096_ & new_n5904_;
  assign new_n5973_ = ~new_n5971_ & ~new_n5972_;
  assign new_n5974_ = lo0040 & new_n5071_;
  assign new_n5975_ = lo0040 & new_n4219_;
  assign new_n5976_ = ~new_n5074_ & new_n5975_;
  assign new_n5977_ = ~new_n5076_ & new_n5956_;
  assign new_n5978_ = ~new_n5976_ & ~new_n5977_;
  assign new_n5979_ = new_n4475_ & ~new_n5978_;
  assign new_n5980_ = lo0040 & new_n5083_;
  assign new_n5981_ = ~new_n5974_ & ~new_n5979_;
  assign new_n5982_ = ~new_n5980_ & new_n5981_;
  assign new_n5983_ = new_n5070_ & ~new_n5982_;
  assign new_n5984_ = ~new_n4096_ & new_n5900_;
  assign new_n5985_ = lo0040 & ~new_n5900_;
  assign new_n5986_ = ~new_n5984_ & ~new_n5985_;
  assign new_n5987_ = new_n5090_ & ~new_n5986_;
  assign new_n5988_ = new_n3746_ & new_n5913_;
  assign new_n5989_ = ~new_n5987_ & ~new_n5988_;
  assign new_n5990_ = new_n5973_ & ~new_n5983_;
  assign new_n5991_ = new_n5989_ & new_n5990_;
  assign new_n5992_ = new_n3804_ & new_n5900_;
  assign new_n5993_ = new_n3834_ & new_n5956_;
  assign new_n5994_ = new_n3678_ & new_n5993_;
  assign new_n5995_ = lo0040 & new_n5112_;
  assign new_n5996_ = new_n3810_ & new_n5904_;
  assign new_n5997_ = ~new_n5992_ & ~new_n5994_;
  assign new_n5998_ = ~new_n5995_ & new_n5997_;
  assign new_n5999_ = ~new_n5996_ & new_n5998_;
  assign new_n6000_ = ~new_n5105_ & new_n5904_;
  assign new_n6001_ = new_n5999_ & ~new_n6000_;
  assign new_n6002_ = new_n3815_ & new_n5913_;
  assign new_n6003_ = new_n4088_ & new_n5900_;
  assign new_n6004_ = ~new_n6002_ & ~new_n6003_;
  assign new_n6005_ = new_n3820_ & new_n5904_;
  assign new_n6006_ = new_n3870_ & new_n5927_;
  assign new_n6007_ = ~new_n6005_ & ~new_n6006_;
  assign new_n6008_ = ~new_n4069_ & new_n5900_;
  assign new_n6009_ = new_n6001_ & new_n6004_;
  assign new_n6010_ = new_n6007_ & new_n6009_;
  assign new_n6011_ = ~new_n6008_ & new_n6010_;
  assign new_n6012_ = new_n5991_ & new_n6011_;
  assign li0040 = ~new_n5970_ | ~new_n6012_;
  assign new_n6014_ = ~new_n4634_ & ~new_n4662_;
  assign new_n6015_ = new_n4642_ & new_n6014_;
  assign new_n6016_ = ~new_n4649_ & new_n6015_;
  assign new_n6017_ = ~new_n4651_ & ~new_n4657_;
  assign new_n6018_ = lo0228 & new_n6017_;
  assign new_n6019_ = ~lo0480 & lo0949;
  assign new_n6020_ = new_n4001_ & new_n6019_;
  assign new_n6021_ = ~lo0250 & lo0252;
  assign new_n6022_ = lo0959 & new_n6021_;
  assign new_n6023_ = new_n3705_ & new_n6022_;
  assign new_n6024_ = lo0901 & new_n6023_;
  assign li0480 = new_n6020_ | new_n6024_;
  assign new_n6026_ = ~lo0228 & ~li0480;
  assign new_n6027_ = new_n6016_ & new_n6018_;
  assign new_n6028_ = ~new_n6026_ & ~new_n6027_;
  assign new_n6029_ = ~lo0044 & ~lo0101;
  assign new_n6030_ = ~lo0041 & new_n6029_;
  assign new_n6031_ = lo0041 & ~new_n6029_;
  assign new_n6032_ = ~new_n6030_ & ~new_n6031_;
  assign new_n6033_ = new_n6028_ & ~new_n6032_;
  assign new_n6034_ = lo0041 & ~new_n6028_;
  assign new_n6035_ = ~new_n6033_ & ~new_n6034_;
  assign new_n6036_ = lo0039 & new_n5253_;
  assign new_n6037_ = new_n3645_ & new_n4543_;
  assign new_n6038_ = ~new_n5323_ & new_n6037_;
  assign new_n6039_ = new_n6036_ & new_n6038_;
  assign new_n6040_ = ~lo0039 & ~new_n6035_;
  assign new_n6041_ = ~new_n6039_ & ~new_n6040_;
  assign li0041 = lo0072 | ~new_n6041_;
  assign new_n6043_ = ~lo0113 & ~lo0116;
  assign new_n6044_ = ~lo0099 & new_n6030_;
  assign new_n6045_ = ~lo0114 & ~lo0115;
  assign new_n6046_ = new_n6043_ & new_n6044_;
  assign new_n6047_ = new_n6045_ & new_n6046_;
  assign new_n6048_ = ~lo0042 & ~new_n6047_;
  assign new_n6049_ = lo0042 & new_n6047_;
  assign new_n6050_ = ~new_n6048_ & ~new_n6049_;
  assign new_n6051_ = lo0042 & ~new_n6028_;
  assign new_n6052_ = new_n6028_ & new_n6050_;
  assign new_n6053_ = ~new_n6051_ & ~new_n6052_;
  assign new_n6054_ = ~lo0039 & ~new_n6053_;
  assign new_n6055_ = lo0200 & new_n3522_;
  assign new_n6056_ = lo0211 & ~new_n3522_;
  assign new_n6057_ = ~new_n6055_ & ~new_n6056_;
  assign new_n6058_ = lo0208 & ~new_n3522_;
  assign new_n6059_ = ~lo0208 & lo0212;
  assign new_n6060_ = ~new_n6058_ & ~new_n6059_;
  assign new_n6061_ = lo0207 & ~new_n3522_;
  assign new_n6062_ = ~lo0207 & lo0214;
  assign new_n6063_ = ~new_n6061_ & ~new_n6062_;
  assign new_n6064_ = new_n6060_ & new_n6063_;
  assign new_n6065_ = ~lo0219 & ~new_n3522_;
  assign new_n6066_ = ~lo0199 & new_n3522_;
  assign new_n6067_ = ~new_n6065_ & ~new_n6066_;
  assign new_n6068_ = ~new_n6057_ & new_n6064_;
  assign new_n6069_ = ~new_n6067_ & ~new_n6068_;
  assign new_n6070_ = lo0039 & ~new_n6037_;
  assign new_n6071_ = ~new_n6069_ & new_n6070_;
  assign new_n6072_ = ~new_n6054_ & ~new_n6071_;
  assign li0042 = ~lo0072 & ~new_n6072_;
  assign new_n6074_ = new_n6057_ & ~new_n6067_;
  assign new_n6075_ = new_n6064_ & new_n6074_;
  assign new_n6076_ = ~new_n6057_ & ~new_n6060_;
  assign new_n6077_ = ~new_n6075_ & ~new_n6076_;
  assign new_n6078_ = ~new_n6037_ & ~new_n6063_;
  assign new_n6079_ = ~new_n6057_ & new_n6078_;
  assign new_n6080_ = ~new_n6037_ & ~new_n6077_;
  assign new_n6081_ = ~new_n6079_ & ~new_n6080_;
  assign new_n6082_ = lo0039 & ~new_n6081_;
  assign new_n6083_ = ~lo0041 & ~lo0101;
  assign new_n6084_ = new_n3657_ & new_n6083_;
  assign new_n6085_ = ~lo0044 & new_n6084_;
  assign new_n6086_ = ~lo0042 & new_n6085_;
  assign new_n6087_ = new_n3656_ & new_n6086_;
  assign new_n6088_ = ~lo0114 & new_n6087_;
  assign new_n6089_ = ~lo0043 & ~new_n6088_;
  assign new_n6090_ = lo0043 & new_n6088_;
  assign new_n6091_ = ~new_n6089_ & ~new_n6090_;
  assign new_n6092_ = lo0043 & ~new_n6028_;
  assign new_n6093_ = new_n6028_ & new_n6091_;
  assign new_n6094_ = ~new_n6092_ & ~new_n6093_;
  assign new_n6095_ = ~lo0039 & ~new_n6094_;
  assign new_n6096_ = ~new_n6082_ & ~new_n6095_;
  assign li0043 = ~lo0072 & ~new_n6096_;
  assign new_n6098_ = lo0044 & ~new_n6028_;
  assign new_n6099_ = ~lo0044 & new_n6028_;
  assign new_n6100_ = ~new_n6098_ & ~new_n6099_;
  assign new_n6101_ = ~lo0039 & ~new_n6100_;
  assign new_n6102_ = new_n5323_ & new_n6037_;
  assign new_n6103_ = new_n6036_ & new_n6102_;
  assign new_n6104_ = ~new_n6101_ & ~new_n6103_;
  assign li0044 = ~lo0072 & ~new_n6104_;
  assign new_n6106_ = lo0045 & ~lo0841;
  assign new_n6107_ = ~lo0024 & lo0045;
  assign new_n6108_ = new_n3804_ & new_n6107_;
  assign new_n6109_ = lo0045 & li0583;
  assign new_n6110_ = new_n3834_ & new_n6109_;
  assign new_n6111_ = new_n3678_ & new_n6110_;
  assign new_n6112_ = lo0045 & new_n5112_;
  assign new_n6113_ = new_n3810_ & new_n6106_;
  assign new_n6114_ = ~new_n6108_ & ~new_n6111_;
  assign new_n6115_ = ~new_n6112_ & new_n6114_;
  assign new_n6116_ = ~new_n6113_ & new_n6115_;
  assign new_n6117_ = ~new_n5105_ & new_n6106_;
  assign new_n6118_ = new_n6116_ & ~new_n6117_;
  assign new_n6119_ = lo0045 & ~lo0314;
  assign new_n6120_ = new_n3815_ & new_n6119_;
  assign new_n6121_ = new_n4088_ & new_n6107_;
  assign new_n6122_ = ~new_n6120_ & ~new_n6121_;
  assign new_n6123_ = ~lo1044 & new_n6119_;
  assign new_n6124_ = new_n3820_ & new_n6106_;
  assign new_n6125_ = new_n3870_ & new_n6123_;
  assign new_n6126_ = ~new_n6124_ & ~new_n6125_;
  assign new_n6127_ = ~new_n4069_ & new_n6107_;
  assign new_n6128_ = new_n6118_ & new_n6122_;
  assign new_n6129_ = new_n6126_ & new_n6128_;
  assign new_n6130_ = ~new_n6127_ & new_n6129_;
  assign new_n6131_ = lo0045 & new_n5194_;
  assign new_n6132_ = ~new_n6107_ & ~new_n6131_;
  assign new_n6133_ = new_n3936_ & ~new_n6132_;
  assign new_n6134_ = new_n3625_ & new_n6107_;
  assign new_n6135_ = ~new_n6133_ & ~new_n6134_;
  assign new_n6136_ = lo0045 & new_n3706_;
  assign new_n6137_ = lo0045 & new_n5608_;
  assign new_n6138_ = ~new_n5184_ & new_n6137_;
  assign new_n6139_ = new_n6135_ & ~new_n6136_;
  assign new_n6140_ = ~new_n6138_ & new_n6139_;
  assign new_n6141_ = ~new_n5201_ & new_n6106_;
  assign new_n6142_ = new_n6140_ & ~new_n6141_;
  assign new_n6143_ = new_n6130_ & new_n6142_;
  assign new_n6144_ = ~new_n5060_ & new_n6119_;
  assign new_n6145_ = new_n3940_ & new_n6107_;
  assign new_n6146_ = ~new_n6144_ & ~new_n6145_;
  assign new_n6147_ = new_n4050_ & new_n6107_;
  assign new_n6148_ = lo0045 & new_n5562_;
  assign new_n6149_ = lo0045 & new_n5155_;
  assign new_n6150_ = new_n3777_ & new_n6149_;
  assign new_n6151_ = lo0045 & ~new_n4632_;
  assign new_n6152_ = new_n5565_ & new_n6151_;
  assign new_n6153_ = ~new_n6150_ & ~new_n6152_;
  assign new_n6154_ = ~new_n5460_ & new_n6119_;
  assign new_n6155_ = new_n6153_ & ~new_n6154_;
  assign new_n6156_ = new_n3763_ & new_n6106_;
  assign new_n6157_ = new_n3780_ & new_n6107_;
  assign new_n6158_ = ~new_n6156_ & ~new_n6157_;
  assign new_n6159_ = new_n3794_ & new_n6119_;
  assign new_n6160_ = new_n6158_ & ~new_n6159_;
  assign new_n6161_ = ~new_n6147_ & ~new_n6148_;
  assign new_n6162_ = new_n6155_ & new_n6161_;
  assign new_n6163_ = new_n6160_ & new_n6162_;
  assign new_n6164_ = new_n4041_ & new_n6107_;
  assign new_n6165_ = new_n6163_ & ~new_n6164_;
  assign new_n6166_ = lo0045 & ~new_n5216_;
  assign new_n6167_ = new_n4133_ & new_n6107_;
  assign new_n6168_ = ~new_n6166_ & ~new_n6167_;
  assign new_n6169_ = new_n3974_ & new_n6109_;
  assign new_n6170_ = ~new_n4135_ & new_n6169_;
  assign new_n6171_ = lo0045 & new_n5225_;
  assign new_n6172_ = new_n6168_ & ~new_n6170_;
  assign new_n6173_ = ~new_n6171_ & new_n6172_;
  assign new_n6174_ = new_n3948_ & new_n6107_;
  assign new_n6175_ = new_n6173_ & ~new_n6174_;
  assign new_n6176_ = lo0045 & new_n3678_;
  assign new_n6177_ = new_n3786_ & new_n6107_;
  assign new_n6178_ = new_n5139_ & new_n6176_;
  assign new_n6179_ = ~new_n6177_ & ~new_n6178_;
  assign new_n6180_ = new_n6146_ & new_n6165_;
  assign new_n6181_ = new_n6175_ & new_n6180_;
  assign new_n6182_ = new_n6179_ & new_n6181_;
  assign new_n6183_ = lo0045 & new_n5135_;
  assign new_n6184_ = new_n4007_ & new_n6123_;
  assign new_n6185_ = new_n3969_ & new_n6106_;
  assign new_n6186_ = ~new_n6184_ & ~new_n6185_;
  assign new_n6187_ = ~new_n6183_ & new_n6186_;
  assign new_n6188_ = lo0045 & new_n5505_;
  assign new_n6189_ = lo0045 & ~lo0993;
  assign new_n6190_ = new_n3927_ & new_n6189_;
  assign new_n6191_ = new_n3953_ & new_n6107_;
  assign new_n6192_ = ~new_n6190_ & ~new_n6191_;
  assign new_n6193_ = new_n6187_ & ~new_n6188_;
  assign new_n6194_ = new_n6192_ & new_n6193_;
  assign new_n6195_ = new_n4020_ & new_n6107_;
  assign new_n6196_ = ~new_n5096_ & new_n6106_;
  assign new_n6197_ = ~new_n6195_ & ~new_n6196_;
  assign new_n6198_ = ~new_n4096_ & new_n6107_;
  assign new_n6199_ = lo0045 & ~new_n6107_;
  assign new_n6200_ = ~new_n6198_ & ~new_n6199_;
  assign new_n6201_ = new_n5090_ & ~new_n6200_;
  assign new_n6202_ = lo0045 & new_n5071_;
  assign new_n6203_ = lo0045 & new_n4219_;
  assign new_n6204_ = ~new_n5074_ & new_n6203_;
  assign new_n6205_ = ~new_n5076_ & new_n6109_;
  assign new_n6206_ = ~new_n6204_ & ~new_n6205_;
  assign new_n6207_ = new_n4475_ & ~new_n6206_;
  assign new_n6208_ = lo0045 & new_n5083_;
  assign new_n6209_ = ~new_n6202_ & ~new_n6207_;
  assign new_n6210_ = ~new_n6208_ & new_n6209_;
  assign new_n6211_ = new_n3612_ & ~new_n6210_;
  assign new_n6212_ = new_n4526_ & new_n6211_;
  assign new_n6213_ = ~lo0287 & new_n6212_;
  assign new_n6214_ = ~lo0287 & lo0979;
  assign new_n6215_ = new_n3612_ & new_n6214_;
  assign new_n6216_ = new_n3746_ & new_n6119_;
  assign new_n6217_ = ~new_n6215_ & ~new_n6216_;
  assign new_n6218_ = new_n6197_ & ~new_n6201_;
  assign new_n6219_ = ~new_n6213_ & new_n6218_;
  assign new_n6220_ = new_n6217_ & new_n6219_;
  assign new_n6221_ = new_n6194_ & new_n6220_;
  assign new_n6222_ = new_n6143_ & new_n6182_;
  assign li0045 = ~new_n6221_ | ~new_n6222_;
  assign new_n6224_ = lo0046 & ~lo0841;
  assign new_n6225_ = ~lo0024 & lo0046;
  assign new_n6226_ = new_n3804_ & new_n6225_;
  assign new_n6227_ = lo0046 & li0583;
  assign new_n6228_ = new_n3834_ & new_n6227_;
  assign new_n6229_ = new_n3678_ & new_n6228_;
  assign new_n6230_ = lo0046 & new_n5112_;
  assign new_n6231_ = new_n3810_ & new_n6224_;
  assign new_n6232_ = ~new_n6226_ & ~new_n6229_;
  assign new_n6233_ = ~new_n6230_ & new_n6232_;
  assign new_n6234_ = ~new_n6231_ & new_n6233_;
  assign new_n6235_ = ~new_n5105_ & new_n6224_;
  assign new_n6236_ = new_n6234_ & ~new_n6235_;
  assign new_n6237_ = lo0046 & ~lo0314;
  assign new_n6238_ = new_n3815_ & new_n6237_;
  assign new_n6239_ = new_n4088_ & new_n6225_;
  assign new_n6240_ = ~new_n6238_ & ~new_n6239_;
  assign new_n6241_ = ~lo1044 & new_n6237_;
  assign new_n6242_ = new_n3820_ & new_n6224_;
  assign new_n6243_ = new_n3870_ & new_n6241_;
  assign new_n6244_ = ~new_n6242_ & ~new_n6243_;
  assign new_n6245_ = ~new_n4069_ & new_n6225_;
  assign new_n6246_ = new_n6236_ & new_n6240_;
  assign new_n6247_ = new_n6244_ & new_n6246_;
  assign new_n6248_ = ~new_n6245_ & new_n6247_;
  assign new_n6249_ = lo0046 & new_n5194_;
  assign new_n6250_ = ~new_n6225_ & ~new_n6249_;
  assign new_n6251_ = new_n3936_ & ~new_n6250_;
  assign new_n6252_ = new_n3625_ & new_n6225_;
  assign new_n6253_ = ~new_n6251_ & ~new_n6252_;
  assign new_n6254_ = lo0046 & new_n3706_;
  assign new_n6255_ = lo0046 & new_n5608_;
  assign new_n6256_ = ~new_n5184_ & new_n6255_;
  assign new_n6257_ = new_n6253_ & ~new_n6254_;
  assign new_n6258_ = ~new_n6256_ & new_n6257_;
  assign new_n6259_ = ~new_n5201_ & new_n6224_;
  assign new_n6260_ = new_n6258_ & ~new_n6259_;
  assign new_n6261_ = new_n6248_ & new_n6260_;
  assign new_n6262_ = lo0046 & new_n5135_;
  assign new_n6263_ = new_n4007_ & new_n6241_;
  assign new_n6264_ = new_n3969_ & new_n6224_;
  assign new_n6265_ = ~new_n6263_ & ~new_n6264_;
  assign new_n6266_ = ~new_n6262_ & new_n6265_;
  assign new_n6267_ = lo0046 & new_n5505_;
  assign new_n6268_ = lo0046 & ~lo0993;
  assign new_n6269_ = new_n3927_ & new_n6268_;
  assign new_n6270_ = new_n3953_ & new_n6225_;
  assign new_n6271_ = ~new_n6269_ & ~new_n6270_;
  assign new_n6272_ = new_n6266_ & ~new_n6267_;
  assign new_n6273_ = new_n6271_ & new_n6272_;
  assign new_n6274_ = lo0046 & new_n5071_;
  assign new_n6275_ = lo0046 & new_n4219_;
  assign new_n6276_ = ~new_n5074_ & new_n6275_;
  assign new_n6277_ = ~new_n5076_ & new_n6227_;
  assign new_n6278_ = ~new_n6276_ & ~new_n6277_;
  assign new_n6279_ = new_n4475_ & ~new_n6278_;
  assign new_n6280_ = lo0046 & new_n5083_;
  assign new_n6281_ = ~new_n6274_ & ~new_n6279_;
  assign new_n6282_ = ~new_n6280_ & new_n6281_;
  assign new_n6283_ = new_n5070_ & ~new_n6282_;
  assign new_n6284_ = new_n4096_ & ~new_n6225_;
  assign new_n6285_ = ~lo0046 & ~new_n4096_;
  assign new_n6286_ = ~new_n6284_ & ~new_n6285_;
  assign new_n6287_ = ~lo0046 & ~lo0841;
  assign new_n6288_ = new_n5090_ & new_n6286_;
  assign new_n6289_ = new_n3735_ & ~new_n6287_;
  assign new_n6290_ = ~new_n6288_ & ~new_n6289_;
  assign new_n6291_ = ~new_n6283_ & new_n6290_;
  assign new_n6292_ = new_n3746_ & new_n6237_;
  assign new_n6293_ = new_n6291_ & ~new_n6292_;
  assign new_n6294_ = new_n4020_ & new_n6225_;
  assign new_n6295_ = new_n3589_ & new_n6224_;
  assign new_n6296_ = new_n6293_ & ~new_n6294_;
  assign new_n6297_ = ~new_n6295_ & new_n6296_;
  assign new_n6298_ = new_n6273_ & new_n6297_;
  assign new_n6299_ = ~new_n5060_ & new_n6237_;
  assign new_n6300_ = new_n3940_ & new_n6225_;
  assign new_n6301_ = ~new_n6299_ & ~new_n6300_;
  assign new_n6302_ = new_n4050_ & new_n6225_;
  assign new_n6303_ = lo0046 & new_n5562_;
  assign new_n6304_ = lo0046 & new_n5155_;
  assign new_n6305_ = new_n3777_ & new_n6304_;
  assign new_n6306_ = lo0046 & ~new_n4632_;
  assign new_n6307_ = new_n5565_ & new_n6306_;
  assign new_n6308_ = ~new_n6305_ & ~new_n6307_;
  assign new_n6309_ = ~new_n5460_ & new_n6237_;
  assign new_n6310_ = new_n6308_ & ~new_n6309_;
  assign new_n6311_ = new_n3763_ & new_n6224_;
  assign new_n6312_ = new_n3780_ & new_n6225_;
  assign new_n6313_ = ~new_n6311_ & ~new_n6312_;
  assign new_n6314_ = new_n3794_ & new_n6237_;
  assign new_n6315_ = new_n6313_ & ~new_n6314_;
  assign new_n6316_ = ~new_n6302_ & ~new_n6303_;
  assign new_n6317_ = new_n6310_ & new_n6316_;
  assign new_n6318_ = new_n6315_ & new_n6317_;
  assign new_n6319_ = new_n4041_ & new_n6225_;
  assign new_n6320_ = new_n6318_ & ~new_n6319_;
  assign new_n6321_ = lo0046 & ~new_n5216_;
  assign new_n6322_ = new_n4133_ & new_n6225_;
  assign new_n6323_ = ~new_n6321_ & ~new_n6322_;
  assign new_n6324_ = new_n3974_ & new_n6227_;
  assign new_n6325_ = ~new_n4135_ & new_n6324_;
  assign new_n6326_ = lo0046 & new_n5225_;
  assign new_n6327_ = new_n6323_ & ~new_n6325_;
  assign new_n6328_ = ~new_n6326_ & new_n6327_;
  assign new_n6329_ = new_n3948_ & new_n6225_;
  assign new_n6330_ = new_n6328_ & ~new_n6329_;
  assign new_n6331_ = lo0046 & new_n3678_;
  assign new_n6332_ = new_n3786_ & new_n6225_;
  assign new_n6333_ = new_n5139_ & new_n6331_;
  assign new_n6334_ = ~new_n6332_ & ~new_n6333_;
  assign new_n6335_ = new_n6301_ & new_n6320_;
  assign new_n6336_ = new_n6330_ & new_n6335_;
  assign new_n6337_ = new_n6334_ & new_n6336_;
  assign new_n6338_ = new_n6261_ & new_n6298_;
  assign li0046 = ~new_n6337_ | ~new_n6338_;
  assign new_n6340_ = lo0047 & ~lo0841;
  assign new_n6341_ = lo0047 & ~lo0314;
  assign new_n6342_ = new_n3746_ & new_n6341_;
  assign new_n6343_ = ~lo0024 & lo0047;
  assign new_n6344_ = new_n4020_ & new_n6343_;
  assign new_n6345_ = ~new_n6342_ & ~new_n6344_;
  assign new_n6346_ = ~new_n5096_ & new_n6340_;
  assign new_n6347_ = new_n6345_ & ~new_n6346_;
  assign new_n6348_ = lo0047 & li0583;
  assign new_n6349_ = new_n3678_ & ~new_n6348_;
  assign new_n6350_ = new_n3834_ & ~new_n6349_;
  assign new_n6351_ = new_n3804_ & new_n6343_;
  assign new_n6352_ = ~new_n6350_ & ~new_n6351_;
  assign new_n6353_ = new_n3810_ & new_n6340_;
  assign new_n6354_ = lo0047 & new_n5112_;
  assign new_n6355_ = new_n6352_ & ~new_n6353_;
  assign new_n6356_ = ~new_n6354_ & new_n6355_;
  assign new_n6357_ = ~new_n5105_ & new_n6340_;
  assign new_n6358_ = new_n6356_ & ~new_n6357_;
  assign new_n6359_ = new_n3815_ & new_n6341_;
  assign new_n6360_ = new_n4088_ & new_n6343_;
  assign new_n6361_ = ~new_n6359_ & ~new_n6360_;
  assign new_n6362_ = ~lo1044 & new_n6341_;
  assign new_n6363_ = new_n3820_ & new_n6340_;
  assign new_n6364_ = new_n3870_ & new_n6362_;
  assign new_n6365_ = ~new_n6363_ & ~new_n6364_;
  assign new_n6366_ = ~new_n4069_ & new_n6343_;
  assign new_n6367_ = new_n6365_ & ~new_n6366_;
  assign new_n6368_ = new_n6347_ & new_n6358_;
  assign new_n6369_ = new_n6361_ & new_n6368_;
  assign new_n6370_ = new_n6367_ & new_n6369_;
  assign new_n6371_ = lo0047 & new_n5071_;
  assign new_n6372_ = lo0047 & lo0786;
  assign new_n6373_ = ~new_n5076_ & new_n6348_;
  assign new_n6374_ = lo0047 & new_n5545_;
  assign new_n6375_ = ~new_n6373_ & ~new_n6374_;
  assign new_n6376_ = new_n4475_ & ~new_n6375_;
  assign new_n6377_ = new_n5082_ & new_n6372_;
  assign new_n6378_ = ~new_n6376_ & ~new_n6377_;
  assign new_n6379_ = ~new_n6371_ & new_n6378_;
  assign new_n6380_ = new_n5070_ & ~new_n6379_;
  assign new_n6381_ = new_n3753_ & new_n4528_;
  assign new_n6382_ = ~new_n4096_ & new_n6343_;
  assign new_n6383_ = lo0047 & ~new_n6343_;
  assign new_n6384_ = ~new_n6382_ & ~new_n6383_;
  assign new_n6385_ = new_n5090_ & ~new_n6384_;
  assign new_n6386_ = ~new_n6381_ & ~new_n6385_;
  assign new_n6387_ = ~new_n6380_ & new_n6386_;
  assign new_n6388_ = new_n6370_ & new_n6387_;
  assign new_n6389_ = ~new_n3786_ & ~new_n4041_;
  assign new_n6390_ = ~new_n4050_ & new_n6389_;
  assign new_n6391_ = lo0047 & new_n5155_;
  assign new_n6392_ = new_n3777_ & new_n6391_;
  assign new_n6393_ = lo0047 & ~new_n4632_;
  assign new_n6394_ = new_n5565_ & new_n6393_;
  assign new_n6395_ = ~new_n6392_ & ~new_n6394_;
  assign new_n6396_ = ~new_n5460_ & new_n6341_;
  assign new_n6397_ = new_n6395_ & ~new_n6396_;
  assign new_n6398_ = lo0047 & new_n5562_;
  assign new_n6399_ = ~new_n3678_ & ~new_n5137_;
  assign new_n6400_ = lo0047 & ~new_n5137_;
  assign new_n6401_ = ~new_n6399_ & ~new_n6400_;
  assign new_n6402_ = new_n3891_ & ~new_n6401_;
  assign new_n6403_ = new_n3763_ & new_n6340_;
  assign new_n6404_ = new_n3780_ & new_n6343_;
  assign new_n6405_ = ~new_n6403_ & ~new_n6404_;
  assign new_n6406_ = new_n3794_ & new_n6341_;
  assign new_n6407_ = new_n6405_ & ~new_n6406_;
  assign new_n6408_ = new_n6397_ & ~new_n6398_;
  assign new_n6409_ = ~new_n6402_ & new_n6408_;
  assign new_n6410_ = new_n6407_ & new_n6409_;
  assign new_n6411_ = new_n6343_ & ~new_n6390_;
  assign new_n6412_ = new_n6410_ & ~new_n6411_;
  assign new_n6413_ = lo0047 & ~new_n5216_;
  assign new_n6414_ = new_n4133_ & new_n6343_;
  assign new_n6415_ = ~new_n6413_ & ~new_n6414_;
  assign new_n6416_ = new_n3974_ & new_n6348_;
  assign new_n6417_ = ~new_n4135_ & new_n6416_;
  assign new_n6418_ = lo0047 & new_n5225_;
  assign new_n6419_ = new_n6415_ & ~new_n6417_;
  assign new_n6420_ = ~new_n6418_ & new_n6419_;
  assign new_n6421_ = new_n3948_ & new_n6343_;
  assign new_n6422_ = new_n6420_ & ~new_n6421_;
  assign new_n6423_ = new_n4007_ & new_n6362_;
  assign new_n6424_ = new_n3969_ & new_n6340_;
  assign new_n6425_ = ~new_n6423_ & ~new_n6424_;
  assign new_n6426_ = new_n6412_ & new_n6422_;
  assign new_n6427_ = new_n6425_ & new_n6426_;
  assign new_n6428_ = lo0047 & new_n5505_;
  assign new_n6429_ = lo0047 & new_n5135_;
  assign new_n6430_ = lo0047 & new_n5608_;
  assign new_n6431_ = ~new_n5184_ & new_n6430_;
  assign new_n6432_ = lo0047 & ~li0583;
  assign new_n6433_ = ~new_n4528_ & ~new_n6432_;
  assign new_n6434_ = new_n4631_ & ~new_n6433_;
  assign new_n6435_ = new_n3936_ & new_n6343_;
  assign new_n6436_ = ~new_n6434_ & ~new_n6435_;
  assign new_n6437_ = new_n3625_ & new_n6343_;
  assign new_n6438_ = lo0047 & new_n3706_;
  assign new_n6439_ = ~new_n6431_ & new_n6436_;
  assign new_n6440_ = ~new_n6437_ & new_n6439_;
  assign new_n6441_ = ~new_n6438_ & new_n6440_;
  assign new_n6442_ = ~new_n5201_ & new_n6340_;
  assign new_n6443_ = new_n6441_ & ~new_n6442_;
  assign new_n6444_ = ~new_n6428_ & ~new_n6429_;
  assign new_n6445_ = new_n6443_ & new_n6444_;
  assign new_n6446_ = new_n6427_ & new_n6445_;
  assign new_n6447_ = ~new_n5060_ & new_n6341_;
  assign new_n6448_ = new_n3940_ & new_n6343_;
  assign new_n6449_ = ~new_n6447_ & ~new_n6448_;
  assign new_n6450_ = lo0047 & ~lo0993;
  assign new_n6451_ = new_n3927_ & new_n6450_;
  assign new_n6452_ = new_n3953_ & new_n6343_;
  assign new_n6453_ = ~new_n6451_ & ~new_n6452_;
  assign new_n6454_ = new_n6449_ & new_n6453_;
  assign new_n6455_ = new_n6388_ & new_n6446_;
  assign li0047 = ~new_n6454_ | ~new_n6455_;
  assign new_n6457_ = lo0048 & new_n5135_;
  assign new_n6458_ = lo0048 & ~lo0841;
  assign new_n6459_ = lo0048 & ~lo0314;
  assign new_n6460_ = ~lo1044 & new_n6459_;
  assign new_n6461_ = new_n4007_ & new_n6460_;
  assign new_n6462_ = new_n3969_ & new_n6458_;
  assign new_n6463_ = ~new_n6461_ & ~new_n6462_;
  assign new_n6464_ = ~new_n6457_ & new_n6463_;
  assign new_n6465_ = lo0048 & new_n5505_;
  assign new_n6466_ = lo0048 & ~lo0993;
  assign new_n6467_ = ~lo0024 & lo0048;
  assign new_n6468_ = new_n3927_ & new_n6466_;
  assign new_n6469_ = new_n3953_ & new_n6467_;
  assign new_n6470_ = ~new_n6468_ & ~new_n6469_;
  assign new_n6471_ = new_n6464_ & ~new_n6465_;
  assign new_n6472_ = new_n6470_ & new_n6471_;
  assign new_n6473_ = new_n4020_ & new_n6467_;
  assign new_n6474_ = ~new_n5096_ & new_n6458_;
  assign new_n6475_ = ~new_n6473_ & ~new_n6474_;
  assign new_n6476_ = lo0048 & new_n5071_;
  assign new_n6477_ = lo0048 & new_n4219_;
  assign new_n6478_ = lo0048 & li0583;
  assign new_n6479_ = ~new_n5074_ & new_n6477_;
  assign new_n6480_ = ~new_n5076_ & new_n6478_;
  assign new_n6481_ = ~new_n6479_ & ~new_n6480_;
  assign new_n6482_ = new_n4475_ & ~new_n6481_;
  assign new_n6483_ = lo0048 & new_n5083_;
  assign new_n6484_ = ~new_n6476_ & ~new_n6482_;
  assign new_n6485_ = ~new_n6483_ & new_n6484_;
  assign new_n6486_ = new_n5070_ & ~new_n6485_;
  assign new_n6487_ = ~new_n4096_ & new_n6467_;
  assign new_n6488_ = lo0048 & ~new_n6467_;
  assign new_n6489_ = ~new_n6487_ & ~new_n6488_;
  assign new_n6490_ = new_n5090_ & ~new_n6489_;
  assign new_n6491_ = new_n3746_ & new_n6459_;
  assign new_n6492_ = ~new_n6490_ & ~new_n6491_;
  assign new_n6493_ = new_n6475_ & ~new_n6486_;
  assign new_n6494_ = new_n6492_ & new_n6493_;
  assign new_n6495_ = new_n6472_ & new_n6494_;
  assign new_n6496_ = lo0048 & new_n5194_;
  assign new_n6497_ = ~new_n6467_ & ~new_n6496_;
  assign new_n6498_ = new_n3936_ & ~new_n6497_;
  assign new_n6499_ = new_n3625_ & new_n6467_;
  assign new_n6500_ = ~new_n6498_ & ~new_n6499_;
  assign new_n6501_ = lo0048 & new_n3706_;
  assign new_n6502_ = lo0048 & new_n5608_;
  assign new_n6503_ = ~new_n5184_ & new_n6502_;
  assign new_n6504_ = new_n6500_ & ~new_n6501_;
  assign new_n6505_ = ~new_n6503_ & new_n6504_;
  assign new_n6506_ = ~new_n5201_ & new_n6458_;
  assign new_n6507_ = new_n6505_ & ~new_n6506_;
  assign new_n6508_ = ~new_n5060_ & new_n6459_;
  assign new_n6509_ = new_n3940_ & new_n6467_;
  assign new_n6510_ = ~new_n6508_ & ~new_n6509_;
  assign new_n6511_ = new_n6507_ & new_n6510_;
  assign new_n6512_ = new_n4050_ & new_n6467_;
  assign new_n6513_ = lo0048 & new_n5562_;
  assign new_n6514_ = lo0048 & new_n5155_;
  assign new_n6515_ = new_n3777_ & new_n6514_;
  assign new_n6516_ = lo0048 & ~new_n4632_;
  assign new_n6517_ = new_n5565_ & new_n6516_;
  assign new_n6518_ = ~new_n6515_ & ~new_n6517_;
  assign new_n6519_ = ~new_n5460_ & new_n6459_;
  assign new_n6520_ = new_n6518_ & ~new_n6519_;
  assign new_n6521_ = new_n3763_ & new_n6458_;
  assign new_n6522_ = new_n3780_ & new_n6467_;
  assign new_n6523_ = ~new_n6521_ & ~new_n6522_;
  assign new_n6524_ = new_n3794_ & new_n6459_;
  assign new_n6525_ = new_n6523_ & ~new_n6524_;
  assign new_n6526_ = ~new_n6512_ & ~new_n6513_;
  assign new_n6527_ = new_n6520_ & new_n6526_;
  assign new_n6528_ = new_n6525_ & new_n6527_;
  assign new_n6529_ = new_n4041_ & new_n6467_;
  assign new_n6530_ = new_n6528_ & ~new_n6529_;
  assign new_n6531_ = lo0048 & ~new_n5216_;
  assign new_n6532_ = new_n4133_ & new_n6467_;
  assign new_n6533_ = ~new_n6531_ & ~new_n6532_;
  assign new_n6534_ = new_n3974_ & new_n6478_;
  assign new_n6535_ = ~new_n4135_ & new_n6534_;
  assign new_n6536_ = lo0048 & new_n5225_;
  assign new_n6537_ = new_n6533_ & ~new_n6535_;
  assign new_n6538_ = ~new_n6536_ & new_n6537_;
  assign new_n6539_ = new_n3948_ & new_n6467_;
  assign new_n6540_ = new_n6538_ & ~new_n6539_;
  assign new_n6541_ = lo0048 & new_n3678_;
  assign new_n6542_ = new_n3786_ & new_n6467_;
  assign new_n6543_ = new_n5139_ & new_n6541_;
  assign new_n6544_ = ~new_n6542_ & ~new_n6543_;
  assign new_n6545_ = new_n6540_ & new_n6544_;
  assign new_n6546_ = new_n6530_ & new_n6545_;
  assign new_n6547_ = new_n3804_ & new_n6467_;
  assign new_n6548_ = new_n3834_ & new_n6478_;
  assign new_n6549_ = new_n3678_ & new_n6548_;
  assign new_n6550_ = lo0048 & new_n5112_;
  assign new_n6551_ = new_n3810_ & new_n6458_;
  assign new_n6552_ = ~new_n6547_ & ~new_n6549_;
  assign new_n6553_ = ~new_n6550_ & new_n6552_;
  assign new_n6554_ = ~new_n6551_ & new_n6553_;
  assign new_n6555_ = ~new_n5105_ & new_n6458_;
  assign new_n6556_ = new_n6554_ & ~new_n6555_;
  assign new_n6557_ = new_n3815_ & new_n6459_;
  assign new_n6558_ = new_n4088_ & new_n6467_;
  assign new_n6559_ = ~new_n6557_ & ~new_n6558_;
  assign new_n6560_ = new_n3820_ & new_n6458_;
  assign new_n6561_ = new_n3870_ & new_n6460_;
  assign new_n6562_ = ~new_n6560_ & ~new_n6561_;
  assign new_n6563_ = ~new_n4069_ & new_n6467_;
  assign new_n6564_ = new_n6556_ & new_n6559_;
  assign new_n6565_ = new_n6562_ & new_n6564_;
  assign new_n6566_ = ~new_n6563_ & new_n6565_;
  assign new_n6567_ = new_n6546_ & new_n6566_;
  assign new_n6568_ = new_n6495_ & new_n6511_;
  assign li0048 = ~new_n6567_ | ~new_n6568_;
  assign new_n6570_ = lo0049 & ~lo0841;
  assign new_n6571_ = ~lo0024 & lo0049;
  assign new_n6572_ = new_n4020_ & new_n6571_;
  assign new_n6573_ = ~new_n5096_ & new_n6570_;
  assign new_n6574_ = ~new_n6572_ & ~new_n6573_;
  assign new_n6575_ = lo0049 & new_n5071_;
  assign new_n6576_ = lo0049 & new_n4219_;
  assign new_n6577_ = lo0049 & li0583;
  assign new_n6578_ = ~new_n5074_ & new_n6576_;
  assign new_n6579_ = ~new_n5076_ & new_n6577_;
  assign new_n6580_ = ~new_n6578_ & ~new_n6579_;
  assign new_n6581_ = new_n4475_ & ~new_n6580_;
  assign new_n6582_ = lo0049 & new_n5083_;
  assign new_n6583_ = ~new_n6575_ & ~new_n6581_;
  assign new_n6584_ = ~new_n6582_ & new_n6583_;
  assign new_n6585_ = new_n5070_ & ~new_n6584_;
  assign new_n6586_ = ~new_n4096_ & new_n6571_;
  assign new_n6587_ = lo0049 & ~new_n6571_;
  assign new_n6588_ = ~new_n6586_ & ~new_n6587_;
  assign new_n6589_ = lo0049 & ~lo0314;
  assign new_n6590_ = new_n5090_ & ~new_n6588_;
  assign new_n6591_ = new_n3746_ & new_n6589_;
  assign new_n6592_ = ~new_n6590_ & ~new_n6591_;
  assign new_n6593_ = new_n6574_ & ~new_n6585_;
  assign new_n6594_ = new_n6592_ & new_n6593_;
  assign new_n6595_ = lo0049 & new_n5112_;
  assign new_n6596_ = new_n3810_ & new_n6570_;
  assign new_n6597_ = new_n3834_ & new_n6577_;
  assign new_n6598_ = new_n3678_ & new_n6597_;
  assign new_n6599_ = ~lo0024 & ~lo0049;
  assign new_n6600_ = new_n4068_ & ~new_n6599_;
  assign new_n6601_ = ~new_n6595_ & ~new_n6596_;
  assign new_n6602_ = ~new_n6598_ & new_n6601_;
  assign new_n6603_ = ~new_n6600_ & new_n6602_;
  assign new_n6604_ = ~new_n5105_ & new_n6570_;
  assign new_n6605_ = new_n6603_ & ~new_n6604_;
  assign new_n6606_ = new_n3815_ & new_n6589_;
  assign new_n6607_ = new_n4088_ & new_n6571_;
  assign new_n6608_ = ~new_n6606_ & ~new_n6607_;
  assign new_n6609_ = ~lo1044 & new_n6589_;
  assign new_n6610_ = new_n3820_ & new_n6570_;
  assign new_n6611_ = new_n3870_ & new_n6609_;
  assign new_n6612_ = ~new_n6610_ & ~new_n6611_;
  assign new_n6613_ = ~new_n3618_ & ~new_n3804_;
  assign new_n6614_ = new_n6571_ & ~new_n6613_;
  assign new_n6615_ = new_n6605_ & new_n6608_;
  assign new_n6616_ = new_n6612_ & new_n6615_;
  assign new_n6617_ = ~new_n6614_ & new_n6616_;
  assign new_n6618_ = new_n6594_ & new_n6617_;
  assign new_n6619_ = ~new_n5060_ & new_n6589_;
  assign new_n6620_ = new_n3940_ & new_n6571_;
  assign new_n6621_ = ~new_n6619_ & ~new_n6620_;
  assign new_n6622_ = lo0049 & ~lo0993;
  assign new_n6623_ = new_n3927_ & new_n6622_;
  assign new_n6624_ = new_n3953_ & new_n6571_;
  assign new_n6625_ = ~new_n6623_ & ~new_n6624_;
  assign new_n6626_ = new_n6621_ & new_n6625_;
  assign new_n6627_ = lo0049 & new_n5194_;
  assign new_n6628_ = ~new_n6571_ & ~new_n6627_;
  assign new_n6629_ = new_n3936_ & ~new_n6628_;
  assign new_n6630_ = new_n3625_ & new_n6571_;
  assign new_n6631_ = ~new_n6629_ & ~new_n6630_;
  assign new_n6632_ = lo0049 & new_n3706_;
  assign new_n6633_ = lo0049 & new_n5608_;
  assign new_n6634_ = ~new_n5184_ & new_n6633_;
  assign new_n6635_ = new_n6631_ & ~new_n6632_;
  assign new_n6636_ = ~new_n6634_ & new_n6635_;
  assign new_n6637_ = ~new_n5201_ & new_n6570_;
  assign new_n6638_ = new_n6636_ & ~new_n6637_;
  assign new_n6639_ = new_n4050_ & new_n6571_;
  assign new_n6640_ = lo0049 & new_n5562_;
  assign new_n6641_ = ~new_n4632_ & new_n5565_;
  assign new_n6642_ = lo0049 & new_n6641_;
  assign new_n6643_ = new_n3777_ & new_n5155_;
  assign new_n6644_ = lo0049 & new_n6643_;
  assign new_n6645_ = ~new_n6642_ & ~new_n6644_;
  assign new_n6646_ = ~new_n5460_ & new_n6589_;
  assign new_n6647_ = new_n6645_ & ~new_n6646_;
  assign new_n6648_ = new_n3763_ & new_n6570_;
  assign new_n6649_ = new_n3780_ & new_n6571_;
  assign new_n6650_ = ~new_n6648_ & ~new_n6649_;
  assign new_n6651_ = new_n3794_ & new_n6589_;
  assign new_n6652_ = new_n6650_ & ~new_n6651_;
  assign new_n6653_ = ~new_n6639_ & ~new_n6640_;
  assign new_n6654_ = new_n6647_ & new_n6653_;
  assign new_n6655_ = new_n6652_ & new_n6654_;
  assign new_n6656_ = new_n4041_ & new_n6571_;
  assign new_n6657_ = new_n6655_ & ~new_n6656_;
  assign new_n6658_ = lo0049 & ~new_n5216_;
  assign new_n6659_ = new_n4133_ & new_n6571_;
  assign new_n6660_ = ~new_n6658_ & ~new_n6659_;
  assign new_n6661_ = new_n3974_ & new_n6577_;
  assign new_n6662_ = ~new_n4135_ & new_n6661_;
  assign new_n6663_ = lo0049 & new_n5225_;
  assign new_n6664_ = new_n6660_ & ~new_n6662_;
  assign new_n6665_ = ~new_n6663_ & new_n6664_;
  assign new_n6666_ = new_n3948_ & new_n6571_;
  assign new_n6667_ = new_n6665_ & ~new_n6666_;
  assign new_n6668_ = lo0049 & new_n3678_;
  assign new_n6669_ = new_n3786_ & new_n6571_;
  assign new_n6670_ = new_n5139_ & new_n6668_;
  assign new_n6671_ = ~new_n6669_ & ~new_n6670_;
  assign new_n6672_ = new_n6657_ & new_n6667_;
  assign new_n6673_ = new_n6671_ & new_n6672_;
  assign new_n6674_ = lo0049 & new_n5505_;
  assign new_n6675_ = lo0049 & new_n5135_;
  assign new_n6676_ = new_n4007_ & new_n6609_;
  assign new_n6677_ = new_n3969_ & new_n6570_;
  assign new_n6678_ = ~new_n6676_ & ~new_n6677_;
  assign new_n6679_ = ~new_n6674_ & ~new_n6675_;
  assign new_n6680_ = new_n6678_ & new_n6679_;
  assign new_n6681_ = new_n6673_ & new_n6680_;
  assign new_n6682_ = new_n6618_ & new_n6626_;
  assign new_n6683_ = new_n6638_ & new_n6682_;
  assign li0049 = ~new_n6681_ | ~new_n6683_;
  assign new_n6685_ = ~new_n3689_ & new_n4647_;
  assign new_n6686_ = ~new_n5182_ & new_n6685_;
  assign new_n6687_ = ~new_n3688_ & ~new_n5184_;
  assign new_n6688_ = lo0050 & new_n6687_;
  assign new_n6689_ = new_n6686_ & new_n6688_;
  assign new_n6690_ = lo0050 & new_n3689_;
  assign new_n6691_ = ~new_n6689_ & ~new_n6690_;
  assign new_n6692_ = ~new_n4581_ & new_n6691_;
  assign new_n6693_ = lo0050 & ~lo0314;
  assign new_n6694_ = ~new_n5060_ & new_n6693_;
  assign new_n6695_ = ~lo0024 & lo0050;
  assign new_n6696_ = new_n3940_ & new_n6695_;
  assign new_n6697_ = ~new_n6694_ & ~new_n6696_;
  assign new_n6698_ = lo0050 & new_n5194_;
  assign new_n6699_ = ~new_n6695_ & ~new_n6698_;
  assign new_n6700_ = new_n3936_ & ~new_n6699_;
  assign new_n6701_ = new_n3625_ & new_n6695_;
  assign new_n6702_ = ~new_n6700_ & ~new_n6701_;
  assign new_n6703_ = lo0050 & ~lo0993;
  assign new_n6704_ = new_n3953_ & new_n6695_;
  assign new_n6705_ = new_n3927_ & new_n6703_;
  assign new_n6706_ = ~new_n6704_ & ~new_n6705_;
  assign new_n6707_ = lo0050 & ~lo0841;
  assign new_n6708_ = ~new_n5201_ & new_n6707_;
  assign new_n6709_ = new_n6697_ & new_n6702_;
  assign new_n6710_ = new_n6706_ & new_n6709_;
  assign new_n6711_ = ~new_n6708_ & new_n6710_;
  assign new_n6712_ = lo0050 & new_n4647_;
  assign new_n6713_ = ~new_n5131_ & ~new_n6712_;
  assign new_n6714_ = ~new_n5134_ & new_n6713_;
  assign new_n6715_ = new_n3705_ & ~new_n6714_;
  assign new_n6716_ = new_n6711_ & ~new_n6715_;
  assign new_n6717_ = new_n3699_ & ~new_n6692_;
  assign new_n6718_ = new_n6716_ & ~new_n6717_;
  assign new_n6719_ = lo0050 & new_n5505_;
  assign new_n6720_ = lo0050 & ~new_n5216_;
  assign new_n6721_ = new_n4133_ & new_n6695_;
  assign new_n6722_ = ~new_n6720_ & ~new_n6721_;
  assign new_n6723_ = lo0050 & li0583;
  assign new_n6724_ = new_n3974_ & new_n6723_;
  assign new_n6725_ = ~new_n4135_ & new_n6724_;
  assign new_n6726_ = lo0050 & new_n5225_;
  assign new_n6727_ = new_n6722_ & ~new_n6725_;
  assign new_n6728_ = ~new_n6726_ & new_n6727_;
  assign new_n6729_ = new_n3948_ & new_n6695_;
  assign new_n6730_ = new_n6728_ & ~new_n6729_;
  assign new_n6731_ = ~lo1044 & new_n6693_;
  assign new_n6732_ = new_n4007_ & new_n6731_;
  assign new_n6733_ = new_n3969_ & new_n6707_;
  assign new_n6734_ = ~new_n6732_ & ~new_n6733_;
  assign new_n6735_ = new_n6730_ & new_n6734_;
  assign new_n6736_ = lo0024 & new_n5170_;
  assign new_n6737_ = ~li0683 & new_n6736_;
  assign new_n6738_ = new_n5171_ & new_n6737_;
  assign new_n6739_ = new_n4050_ & new_n6695_;
  assign new_n6740_ = ~new_n6738_ & ~new_n6739_;
  assign new_n6741_ = lo0050 & new_n5562_;
  assign new_n6742_ = lo0050 & new_n5155_;
  assign new_n6743_ = new_n3777_ & new_n6742_;
  assign new_n6744_ = lo0050 & ~new_n4632_;
  assign new_n6745_ = new_n5565_ & new_n6744_;
  assign new_n6746_ = ~new_n6743_ & ~new_n6745_;
  assign new_n6747_ = ~new_n5460_ & new_n6693_;
  assign new_n6748_ = new_n6746_ & ~new_n6747_;
  assign new_n6749_ = new_n3780_ & new_n6695_;
  assign new_n6750_ = new_n3763_ & new_n6707_;
  assign new_n6751_ = ~new_n6749_ & ~new_n6750_;
  assign new_n6752_ = new_n3794_ & new_n6693_;
  assign new_n6753_ = ~new_n6741_ & new_n6748_;
  assign new_n6754_ = new_n6751_ & new_n6753_;
  assign new_n6755_ = ~new_n6752_ & new_n6754_;
  assign new_n6756_ = new_n6740_ & new_n6755_;
  assign new_n6757_ = lo0050 & new_n5140_;
  assign new_n6758_ = new_n3786_ & new_n6695_;
  assign new_n6759_ = ~new_n6757_ & ~new_n6758_;
  assign new_n6760_ = new_n4041_ & new_n6695_;
  assign new_n6761_ = new_n6759_ & ~new_n6760_;
  assign new_n6762_ = ~new_n6719_ & new_n6735_;
  assign new_n6763_ = new_n6756_ & new_n6762_;
  assign new_n6764_ = new_n6761_ & new_n6763_;
  assign new_n6765_ = new_n6718_ & new_n6764_;
  assign new_n6766_ = new_n3834_ & new_n6723_;
  assign new_n6767_ = new_n3678_ & new_n6766_;
  assign new_n6768_ = new_n3804_ & new_n6695_;
  assign new_n6769_ = ~new_n6767_ & ~new_n6768_;
  assign new_n6770_ = new_n3810_ & new_n6707_;
  assign new_n6771_ = lo0050 & new_n5112_;
  assign new_n6772_ = ~new_n6770_ & ~new_n6771_;
  assign new_n6773_ = new_n6769_ & new_n6772_;
  assign new_n6774_ = new_n4020_ & new_n6695_;
  assign new_n6775_ = ~new_n5096_ & new_n6707_;
  assign new_n6776_ = ~new_n6774_ & ~new_n6775_;
  assign new_n6777_ = ~new_n4096_ & new_n6695_;
  assign new_n6778_ = lo0050 & ~new_n6695_;
  assign new_n6779_ = ~new_n6777_ & ~new_n6778_;
  assign new_n6780_ = new_n5090_ & ~new_n6779_;
  assign new_n6781_ = new_n3746_ & new_n6693_;
  assign new_n6782_ = ~new_n6780_ & ~new_n6781_;
  assign new_n6783_ = lo0050 & new_n5071_;
  assign new_n6784_ = lo0050 & new_n4219_;
  assign new_n6785_ = ~new_n5074_ & new_n6784_;
  assign new_n6786_ = ~new_n5076_ & new_n6723_;
  assign new_n6787_ = ~new_n6785_ & ~new_n6786_;
  assign new_n6788_ = new_n4475_ & ~new_n6787_;
  assign new_n6789_ = lo0050 & new_n5083_;
  assign new_n6790_ = ~new_n6783_ & ~new_n6788_;
  assign new_n6791_ = ~new_n6789_ & new_n6790_;
  assign new_n6792_ = new_n5070_ & ~new_n6791_;
  assign new_n6793_ = new_n6773_ & new_n6776_;
  assign new_n6794_ = new_n6782_ & new_n6793_;
  assign new_n6795_ = ~new_n6792_ & new_n6794_;
  assign new_n6796_ = ~new_n5105_ & new_n6707_;
  assign new_n6797_ = new_n6795_ & ~new_n6796_;
  assign new_n6798_ = new_n3815_ & new_n6693_;
  assign new_n6799_ = new_n4088_ & new_n6695_;
  assign new_n6800_ = ~new_n6798_ & ~new_n6799_;
  assign new_n6801_ = new_n3820_ & new_n6707_;
  assign new_n6802_ = new_n3870_ & new_n6731_;
  assign new_n6803_ = ~new_n6801_ & ~new_n6802_;
  assign new_n6804_ = ~new_n4069_ & new_n6695_;
  assign new_n6805_ = new_n6803_ & ~new_n6804_;
  assign new_n6806_ = new_n6765_ & new_n6797_;
  assign new_n6807_ = new_n6800_ & new_n6806_;
  assign li0050 = ~new_n6805_ | ~new_n6807_;
  assign new_n6809_ = lo0051 & new_n5230_;
  assign new_n6810_ = lo0051 & new_n3678_;
  assign new_n6811_ = ~lo0024 & lo0051;
  assign new_n6812_ = new_n3786_ & new_n6811_;
  assign new_n6813_ = new_n5139_ & new_n6810_;
  assign new_n6814_ = ~new_n6812_ & ~new_n6813_;
  assign new_n6815_ = lo0051 & ~lo0841;
  assign new_n6816_ = lo0051 & ~lo0314;
  assign new_n6817_ = ~lo1044 & new_n6816_;
  assign new_n6818_ = new_n4007_ & new_n6817_;
  assign new_n6819_ = new_n3969_ & new_n6815_;
  assign new_n6820_ = ~new_n6818_ & ~new_n6819_;
  assign new_n6821_ = lo0051 & new_n5135_;
  assign new_n6822_ = new_n6814_ & new_n6820_;
  assign new_n6823_ = ~new_n6821_ & new_n6822_;
  assign new_n6824_ = new_n4001_ & new_n6809_;
  assign new_n6825_ = new_n6823_ & ~new_n6824_;
  assign new_n6826_ = new_n4050_ & new_n6811_;
  assign new_n6827_ = lo0051 & new_n5562_;
  assign new_n6828_ = lo0051 & new_n5155_;
  assign new_n6829_ = new_n3777_ & new_n6828_;
  assign new_n6830_ = lo0051 & ~new_n4632_;
  assign new_n6831_ = new_n5565_ & new_n6830_;
  assign new_n6832_ = ~new_n6829_ & ~new_n6831_;
  assign new_n6833_ = ~new_n5460_ & new_n6816_;
  assign new_n6834_ = new_n6832_ & ~new_n6833_;
  assign new_n6835_ = new_n3763_ & new_n6815_;
  assign new_n6836_ = new_n3780_ & new_n6811_;
  assign new_n6837_ = ~new_n6835_ & ~new_n6836_;
  assign new_n6838_ = new_n3794_ & new_n6816_;
  assign new_n6839_ = new_n6837_ & ~new_n6838_;
  assign new_n6840_ = ~new_n6826_ & ~new_n6827_;
  assign new_n6841_ = new_n6834_ & new_n6840_;
  assign new_n6842_ = new_n6839_ & new_n6841_;
  assign new_n6843_ = new_n4041_ & new_n6811_;
  assign new_n6844_ = new_n6842_ & ~new_n6843_;
  assign new_n6845_ = lo0051 & ~new_n5216_;
  assign new_n6846_ = new_n4133_ & new_n6811_;
  assign new_n6847_ = ~new_n6845_ & ~new_n6846_;
  assign new_n6848_ = lo0051 & li0583;
  assign new_n6849_ = new_n3974_ & new_n6848_;
  assign new_n6850_ = ~new_n4135_ & new_n6849_;
  assign new_n6851_ = lo0051 & new_n5225_;
  assign new_n6852_ = new_n6847_ & ~new_n6850_;
  assign new_n6853_ = ~new_n6851_ & new_n6852_;
  assign new_n6854_ = new_n3948_ & new_n6811_;
  assign new_n6855_ = new_n6853_ & ~new_n6854_;
  assign new_n6856_ = new_n6825_ & new_n6844_;
  assign new_n6857_ = new_n6855_ & new_n6856_;
  assign new_n6858_ = lo0051 & new_n5818_;
  assign new_n6859_ = ~new_n5184_ & new_n6858_;
  assign new_n6860_ = lo0051 & new_n3706_;
  assign new_n6861_ = lo0051 & new_n4135_;
  assign new_n6862_ = lo0024 & new_n6861_;
  assign new_n6863_ = ~new_n6811_ & ~new_n6862_;
  assign new_n6864_ = new_n3936_ & ~new_n6863_;
  assign new_n6865_ = new_n3725_ & new_n6815_;
  assign new_n6866_ = new_n3625_ & new_n6811_;
  assign new_n6867_ = ~new_n6865_ & ~new_n6866_;
  assign new_n6868_ = ~new_n5827_ & new_n6815_;
  assign new_n6869_ = new_n6867_ & ~new_n6868_;
  assign new_n6870_ = ~new_n6860_ & ~new_n6864_;
  assign new_n6871_ = new_n6869_ & new_n6870_;
  assign new_n6872_ = ~new_n3723_ & new_n6871_;
  assign new_n6873_ = ~new_n5060_ & new_n6816_;
  assign new_n6874_ = new_n3940_ & new_n6811_;
  assign new_n6875_ = ~new_n6873_ & ~new_n6874_;
  assign new_n6876_ = new_n3953_ & new_n6811_;
  assign new_n6877_ = lo0051 & new_n5671_;
  assign new_n6878_ = new_n6875_ & ~new_n6876_;
  assign new_n6879_ = ~new_n6877_ & new_n6878_;
  assign new_n6880_ = new_n6872_ & new_n6879_;
  assign new_n6881_ = ~new_n6859_ & new_n6880_;
  assign new_n6882_ = new_n6857_ & new_n6881_;
  assign new_n6883_ = new_n4020_ & new_n6811_;
  assign new_n6884_ = ~new_n5096_ & new_n6815_;
  assign new_n6885_ = ~new_n6883_ & ~new_n6884_;
  assign new_n6886_ = lo0051 & new_n5071_;
  assign new_n6887_ = lo0051 & new_n4219_;
  assign new_n6888_ = ~new_n5074_ & new_n6887_;
  assign new_n6889_ = ~new_n5076_ & new_n6848_;
  assign new_n6890_ = ~new_n6888_ & ~new_n6889_;
  assign new_n6891_ = new_n4475_ & ~new_n6890_;
  assign new_n6892_ = lo0051 & new_n5083_;
  assign new_n6893_ = ~new_n6886_ & ~new_n6891_;
  assign new_n6894_ = ~new_n6892_ & new_n6893_;
  assign new_n6895_ = new_n5070_ & ~new_n6894_;
  assign new_n6896_ = ~new_n4096_ & new_n6811_;
  assign new_n6897_ = lo0051 & ~new_n6811_;
  assign new_n6898_ = ~new_n6896_ & ~new_n6897_;
  assign new_n6899_ = new_n5090_ & ~new_n6898_;
  assign new_n6900_ = new_n3746_ & new_n6816_;
  assign new_n6901_ = ~new_n6899_ & ~new_n6900_;
  assign new_n6902_ = new_n6885_ & ~new_n6895_;
  assign new_n6903_ = new_n6901_ & new_n6902_;
  assign new_n6904_ = new_n3804_ & new_n6811_;
  assign new_n6905_ = new_n3834_ & new_n6848_;
  assign new_n6906_ = new_n3678_ & new_n6905_;
  assign new_n6907_ = lo0051 & new_n5112_;
  assign new_n6908_ = new_n3810_ & new_n6815_;
  assign new_n6909_ = ~new_n6904_ & ~new_n6906_;
  assign new_n6910_ = ~new_n6907_ & new_n6909_;
  assign new_n6911_ = ~new_n6908_ & new_n6910_;
  assign new_n6912_ = ~new_n5105_ & new_n6815_;
  assign new_n6913_ = new_n6911_ & ~new_n6912_;
  assign new_n6914_ = new_n3815_ & new_n6816_;
  assign new_n6915_ = new_n4088_ & new_n6811_;
  assign new_n6916_ = ~new_n6914_ & ~new_n6915_;
  assign new_n6917_ = new_n3820_ & new_n6815_;
  assign new_n6918_ = new_n3870_ & new_n6817_;
  assign new_n6919_ = ~new_n6917_ & ~new_n6918_;
  assign new_n6920_ = ~new_n4069_ & new_n6811_;
  assign new_n6921_ = new_n6913_ & new_n6916_;
  assign new_n6922_ = new_n6919_ & new_n6921_;
  assign new_n6923_ = ~new_n6920_ & new_n6922_;
  assign new_n6924_ = new_n6903_ & new_n6923_;
  assign li0051 = ~new_n6882_ | ~new_n6924_;
  assign new_n6926_ = ~new_n6064_ & new_n6070_;
  assign new_n6927_ = new_n6074_ & new_n6926_;
  assign new_n6928_ = ~lo0116 & new_n3657_;
  assign new_n6929_ = new_n6030_ & new_n6928_;
  assign new_n6930_ = new_n6045_ & new_n6929_;
  assign new_n6931_ = new_n3660_ & new_n6930_;
  assign new_n6932_ = lo0052 & ~new_n6931_;
  assign new_n6933_ = ~lo0052 & new_n6931_;
  assign new_n6934_ = ~new_n6932_ & ~new_n6933_;
  assign new_n6935_ = new_n6028_ & new_n6934_;
  assign new_n6936_ = ~lo0052 & ~new_n6028_;
  assign new_n6937_ = ~lo0039 & ~new_n6935_;
  assign new_n6938_ = ~new_n6936_ & new_n6937_;
  assign new_n6939_ = ~new_n6927_ & ~new_n6938_;
  assign li0052 = ~lo0072 & ~new_n6939_;
  assign new_n6941_ = lo0053 & ~lo0841;
  assign new_n6942_ = ~lo0024 & lo0053;
  assign new_n6943_ = new_n4020_ & new_n6942_;
  assign new_n6944_ = ~new_n5096_ & new_n6941_;
  assign new_n6945_ = ~new_n6943_ & ~new_n6944_;
  assign new_n6946_ = ~new_n4096_ & new_n6942_;
  assign new_n6947_ = lo0053 & ~new_n6942_;
  assign new_n6948_ = ~new_n6946_ & ~new_n6947_;
  assign new_n6949_ = new_n5090_ & ~new_n6948_;
  assign new_n6950_ = ~new_n5071_ & ~new_n5083_;
  assign new_n6951_ = lo0053 & new_n4219_;
  assign new_n6952_ = lo0053 & li0583;
  assign new_n6953_ = ~new_n5074_ & new_n6951_;
  assign new_n6954_ = ~new_n5076_ & new_n6952_;
  assign new_n6955_ = ~new_n6953_ & ~new_n6954_;
  assign new_n6956_ = ~new_n4423_ & new_n4475_;
  assign new_n6957_ = ~new_n6955_ & new_n6956_;
  assign new_n6958_ = ~new_n4423_ & ~new_n6950_;
  assign new_n6959_ = lo0053 & new_n6958_;
  assign new_n6960_ = ~new_n6957_ & ~new_n6959_;
  assign new_n6961_ = new_n4525_ & ~new_n6960_;
  assign new_n6962_ = new_n4421_ & new_n4524_;
  assign new_n6963_ = lo0053 & ~lo0314;
  assign new_n6964_ = new_n3612_ & new_n6962_;
  assign new_n6965_ = new_n3746_ & new_n6963_;
  assign new_n6966_ = ~new_n6964_ & ~new_n6965_;
  assign new_n6967_ = new_n6945_ & ~new_n6949_;
  assign new_n6968_ = ~new_n6961_ & new_n6967_;
  assign new_n6969_ = new_n6966_ & new_n6968_;
  assign new_n6970_ = lo0053 & new_n5194_;
  assign new_n6971_ = ~new_n6942_ & ~new_n6970_;
  assign new_n6972_ = new_n3936_ & ~new_n6971_;
  assign new_n6973_ = new_n3625_ & new_n6942_;
  assign new_n6974_ = ~new_n6972_ & ~new_n6973_;
  assign new_n6975_ = lo0053 & new_n3706_;
  assign new_n6976_ = lo0053 & new_n5818_;
  assign new_n6977_ = ~new_n5184_ & new_n6976_;
  assign new_n6978_ = new_n6974_ & ~new_n6975_;
  assign new_n6979_ = ~new_n6977_ & new_n6978_;
  assign new_n6980_ = ~new_n5201_ & new_n6941_;
  assign new_n6981_ = new_n6979_ & ~new_n6980_;
  assign new_n6982_ = new_n6969_ & new_n6981_;
  assign new_n6983_ = lo0053 & new_n5505_;
  assign new_n6984_ = lo0053 & new_n5135_;
  assign new_n6985_ = lo0053 & ~lo0993;
  assign new_n6986_ = new_n3927_ & new_n6985_;
  assign new_n6987_ = new_n3953_ & new_n6942_;
  assign new_n6988_ = ~new_n6986_ & ~new_n6987_;
  assign new_n6989_ = ~lo1044 & new_n6963_;
  assign new_n6990_ = new_n4007_ & new_n6989_;
  assign new_n6991_ = new_n3969_ & new_n6941_;
  assign new_n6992_ = ~new_n6990_ & ~new_n6991_;
  assign new_n6993_ = ~new_n6983_ & ~new_n6984_;
  assign new_n6994_ = new_n6988_ & new_n6993_;
  assign new_n6995_ = new_n6992_ & new_n6994_;
  assign new_n6996_ = new_n3804_ & new_n6942_;
  assign new_n6997_ = new_n3834_ & new_n6952_;
  assign new_n6998_ = new_n3678_ & new_n6997_;
  assign new_n6999_ = lo0053 & new_n5112_;
  assign new_n7000_ = new_n3810_ & new_n6941_;
  assign new_n7001_ = ~new_n6996_ & ~new_n6998_;
  assign new_n7002_ = ~new_n6999_ & new_n7001_;
  assign new_n7003_ = ~new_n7000_ & new_n7002_;
  assign new_n7004_ = ~new_n5105_ & new_n6941_;
  assign new_n7005_ = new_n7003_ & ~new_n7004_;
  assign new_n7006_ = new_n3815_ & new_n6963_;
  assign new_n7007_ = new_n4088_ & new_n6942_;
  assign new_n7008_ = ~new_n7006_ & ~new_n7007_;
  assign new_n7009_ = new_n3820_ & new_n6941_;
  assign new_n7010_ = new_n3870_ & new_n6989_;
  assign new_n7011_ = ~new_n7009_ & ~new_n7010_;
  assign new_n7012_ = ~new_n4069_ & new_n6942_;
  assign new_n7013_ = new_n7005_ & new_n7008_;
  assign new_n7014_ = new_n7011_ & new_n7013_;
  assign new_n7015_ = ~new_n7012_ & new_n7014_;
  assign new_n7016_ = new_n6995_ & new_n7015_;
  assign new_n7017_ = ~new_n5060_ & new_n6963_;
  assign new_n7018_ = new_n3940_ & new_n6942_;
  assign new_n7019_ = ~new_n7017_ & ~new_n7018_;
  assign new_n7020_ = new_n4050_ & new_n6942_;
  assign new_n7021_ = lo0053 & new_n5562_;
  assign new_n7022_ = lo0053 & new_n5155_;
  assign new_n7023_ = new_n3777_ & new_n7022_;
  assign new_n7024_ = lo0053 & ~new_n4632_;
  assign new_n7025_ = new_n5565_ & new_n7024_;
  assign new_n7026_ = ~new_n7023_ & ~new_n7025_;
  assign new_n7027_ = ~new_n5460_ & new_n6963_;
  assign new_n7028_ = new_n7026_ & ~new_n7027_;
  assign new_n7029_ = new_n3763_ & new_n6941_;
  assign new_n7030_ = new_n3780_ & new_n6942_;
  assign new_n7031_ = ~new_n7029_ & ~new_n7030_;
  assign new_n7032_ = new_n3794_ & new_n6963_;
  assign new_n7033_ = new_n7031_ & ~new_n7032_;
  assign new_n7034_ = ~new_n7020_ & ~new_n7021_;
  assign new_n7035_ = new_n7028_ & new_n7034_;
  assign new_n7036_ = new_n7033_ & new_n7035_;
  assign new_n7037_ = new_n4041_ & new_n6942_;
  assign new_n7038_ = new_n7036_ & ~new_n7037_;
  assign new_n7039_ = lo0053 & ~new_n5216_;
  assign new_n7040_ = new_n4133_ & new_n6942_;
  assign new_n7041_ = ~new_n7039_ & ~new_n7040_;
  assign new_n7042_ = new_n3974_ & new_n6952_;
  assign new_n7043_ = ~new_n4135_ & new_n7042_;
  assign new_n7044_ = lo0053 & new_n5225_;
  assign new_n7045_ = new_n7041_ & ~new_n7043_;
  assign new_n7046_ = ~new_n7044_ & new_n7045_;
  assign new_n7047_ = new_n3948_ & new_n6942_;
  assign new_n7048_ = new_n7046_ & ~new_n7047_;
  assign new_n7049_ = lo0053 & new_n3678_;
  assign new_n7050_ = new_n3786_ & new_n6942_;
  assign new_n7051_ = new_n5139_ & new_n7049_;
  assign new_n7052_ = ~new_n7050_ & ~new_n7051_;
  assign new_n7053_ = new_n7019_ & new_n7038_;
  assign new_n7054_ = new_n7048_ & new_n7053_;
  assign new_n7055_ = new_n7052_ & new_n7054_;
  assign new_n7056_ = new_n6982_ & new_n7016_;
  assign li0053 = ~new_n7055_ | ~new_n7056_;
  assign new_n7058_ = ~lo0024 & lo0054;
  assign new_n7059_ = lo0054 & ~lo0314;
  assign new_n7060_ = lo0054 & new_n5155_;
  assign new_n7061_ = new_n3777_ & new_n7060_;
  assign new_n7062_ = lo0054 & ~new_n4632_;
  assign new_n7063_ = new_n5565_ & new_n7062_;
  assign new_n7064_ = ~new_n7061_ & ~new_n7063_;
  assign new_n7065_ = ~new_n5460_ & new_n7059_;
  assign new_n7066_ = new_n7064_ & ~new_n7065_;
  assign new_n7067_ = lo0054 & new_n5562_;
  assign new_n7068_ = new_n4050_ & new_n7058_;
  assign new_n7069_ = lo0054 & ~lo0841;
  assign new_n7070_ = new_n3763_ & new_n7069_;
  assign new_n7071_ = new_n3780_ & new_n7058_;
  assign new_n7072_ = ~new_n7070_ & ~new_n7071_;
  assign new_n7073_ = new_n3794_ & new_n7059_;
  assign new_n7074_ = new_n7072_ & ~new_n7073_;
  assign new_n7075_ = new_n7066_ & ~new_n7067_;
  assign new_n7076_ = ~new_n7068_ & new_n7075_;
  assign new_n7077_ = new_n7074_ & new_n7076_;
  assign new_n7078_ = new_n4041_ & new_n7058_;
  assign new_n7079_ = new_n7077_ & ~new_n7078_;
  assign new_n7080_ = lo0054 & ~new_n5216_;
  assign new_n7081_ = ~lo0054 & ~lo0841;
  assign new_n7082_ = new_n3969_ & ~new_n7081_;
  assign new_n7083_ = lo0054 & new_n5225_;
  assign new_n7084_ = lo0054 & li0583;
  assign new_n7085_ = new_n3974_ & new_n7084_;
  assign new_n7086_ = ~new_n4135_ & new_n7085_;
  assign new_n7087_ = ~new_n7080_ & ~new_n7082_;
  assign new_n7088_ = ~new_n7083_ & new_n7087_;
  assign new_n7089_ = ~new_n7086_ & new_n7088_;
  assign new_n7090_ = new_n4133_ & new_n7058_;
  assign new_n7091_ = new_n7089_ & ~new_n7090_;
  assign new_n7092_ = lo0054 & new_n3678_;
  assign new_n7093_ = new_n3786_ & new_n7058_;
  assign new_n7094_ = new_n5139_ & new_n7092_;
  assign new_n7095_ = ~new_n7093_ & ~new_n7094_;
  assign new_n7096_ = new_n7079_ & new_n7091_;
  assign new_n7097_ = new_n7095_ & new_n7096_;
  assign new_n7098_ = ~new_n5060_ & new_n7059_;
  assign new_n7099_ = new_n3940_ & new_n7058_;
  assign new_n7100_ = ~new_n7098_ & ~new_n7099_;
  assign new_n7101_ = lo0054 & ~lo0993;
  assign new_n7102_ = new_n3927_ & new_n7101_;
  assign new_n7103_ = new_n3953_ & new_n7058_;
  assign new_n7104_ = ~new_n7102_ & ~new_n7103_;
  assign new_n7105_ = new_n7100_ & new_n7104_;
  assign new_n7106_ = new_n7097_ & new_n7105_;
  assign new_n7107_ = new_n4020_ & new_n7058_;
  assign new_n7108_ = ~new_n5096_ & new_n7069_;
  assign new_n7109_ = ~new_n7107_ & ~new_n7108_;
  assign new_n7110_ = lo0054 & new_n5071_;
  assign new_n7111_ = lo0054 & new_n4219_;
  assign new_n7112_ = ~new_n5074_ & new_n7111_;
  assign new_n7113_ = ~new_n5076_ & new_n7084_;
  assign new_n7114_ = ~new_n7112_ & ~new_n7113_;
  assign new_n7115_ = new_n4475_ & ~new_n7114_;
  assign new_n7116_ = lo0054 & new_n5083_;
  assign new_n7117_ = ~new_n7110_ & ~new_n7115_;
  assign new_n7118_ = ~new_n7116_ & new_n7117_;
  assign new_n7119_ = new_n5070_ & ~new_n7118_;
  assign new_n7120_ = ~new_n4096_ & new_n7058_;
  assign new_n7121_ = lo0054 & ~new_n7058_;
  assign new_n7122_ = ~new_n7120_ & ~new_n7121_;
  assign new_n7123_ = new_n5090_ & ~new_n7122_;
  assign new_n7124_ = new_n3746_ & new_n7059_;
  assign new_n7125_ = ~new_n7123_ & ~new_n7124_;
  assign new_n7126_ = new_n7109_ & ~new_n7119_;
  assign new_n7127_ = new_n7125_ & new_n7126_;
  assign new_n7128_ = lo0054 & new_n5505_;
  assign new_n7129_ = lo0054 & new_n5135_;
  assign new_n7130_ = ~lo1044 & new_n7059_;
  assign new_n7131_ = new_n4007_ & new_n7130_;
  assign new_n7132_ = new_n3948_ & new_n7058_;
  assign new_n7133_ = ~new_n7131_ & ~new_n7132_;
  assign new_n7134_ = ~new_n7128_ & ~new_n7129_;
  assign new_n7135_ = new_n7133_ & new_n7134_;
  assign new_n7136_ = new_n3804_ & new_n7058_;
  assign new_n7137_ = new_n3834_ & new_n7084_;
  assign new_n7138_ = new_n3678_ & new_n7137_;
  assign new_n7139_ = lo0054 & new_n5112_;
  assign new_n7140_ = new_n3810_ & new_n7069_;
  assign new_n7141_ = ~new_n7136_ & ~new_n7138_;
  assign new_n7142_ = ~new_n7139_ & new_n7141_;
  assign new_n7143_ = ~new_n7140_ & new_n7142_;
  assign new_n7144_ = ~new_n5105_ & new_n7069_;
  assign new_n7145_ = new_n7143_ & ~new_n7144_;
  assign new_n7146_ = new_n3815_ & new_n7059_;
  assign new_n7147_ = new_n4088_ & new_n7058_;
  assign new_n7148_ = ~new_n7146_ & ~new_n7147_;
  assign new_n7149_ = new_n3820_ & new_n7069_;
  assign new_n7150_ = new_n3870_ & new_n7130_;
  assign new_n7151_ = ~new_n7149_ & ~new_n7150_;
  assign new_n7152_ = ~new_n4069_ & new_n7058_;
  assign new_n7153_ = new_n7145_ & new_n7148_;
  assign new_n7154_ = new_n7151_ & new_n7153_;
  assign new_n7155_ = ~new_n7152_ & new_n7154_;
  assign new_n7156_ = new_n7135_ & new_n7155_;
  assign new_n7157_ = lo0054 & new_n5194_;
  assign new_n7158_ = ~new_n7058_ & ~new_n7157_;
  assign new_n7159_ = new_n3936_ & ~new_n7158_;
  assign new_n7160_ = new_n3625_ & new_n7058_;
  assign new_n7161_ = ~new_n7159_ & ~new_n7160_;
  assign new_n7162_ = lo0054 & new_n3706_;
  assign new_n7163_ = ~new_n5184_ & new_n5818_;
  assign new_n7164_ = lo0054 & new_n7163_;
  assign new_n7165_ = new_n7161_ & ~new_n7162_;
  assign new_n7166_ = ~new_n7164_ & new_n7165_;
  assign new_n7167_ = ~new_n5201_ & new_n7069_;
  assign new_n7168_ = new_n7166_ & ~new_n7167_;
  assign new_n7169_ = new_n7106_ & new_n7127_;
  assign new_n7170_ = new_n7156_ & new_n7169_;
  assign li0054 = ~new_n7168_ | ~new_n7170_;
  assign new_n7172_ = lo0055 & ~lo0314;
  assign new_n7173_ = ~lo0024 & lo0055;
  assign new_n7174_ = ~new_n5060_ & new_n7172_;
  assign new_n7175_ = new_n3940_ & new_n7173_;
  assign new_n7176_ = ~new_n7174_ & ~new_n7175_;
  assign new_n7177_ = lo0055 & ~lo0841;
  assign new_n7178_ = lo0055 & new_n5194_;
  assign new_n7179_ = ~new_n7173_ & ~new_n7178_;
  assign new_n7180_ = new_n3936_ & ~new_n7179_;
  assign new_n7181_ = new_n3625_ & new_n7173_;
  assign new_n7182_ = ~new_n7180_ & ~new_n7181_;
  assign new_n7183_ = lo0055 & new_n3706_;
  assign new_n7184_ = lo0055 & new_n5818_;
  assign new_n7185_ = ~new_n5184_ & new_n7184_;
  assign new_n7186_ = new_n7182_ & ~new_n7183_;
  assign new_n7187_ = ~new_n7185_ & new_n7186_;
  assign new_n7188_ = ~new_n5201_ & new_n7177_;
  assign new_n7189_ = new_n7187_ & ~new_n7188_;
  assign new_n7190_ = new_n7176_ & new_n7189_;
  assign new_n7191_ = new_n4020_ & new_n7173_;
  assign new_n7192_ = ~new_n5096_ & new_n7177_;
  assign new_n7193_ = ~new_n7191_ & ~new_n7192_;
  assign new_n7194_ = lo0055 & new_n5071_;
  assign new_n7195_ = lo0055 & new_n4219_;
  assign new_n7196_ = lo0055 & li0583;
  assign new_n7197_ = ~new_n5074_ & new_n7195_;
  assign new_n7198_ = ~new_n5076_ & new_n7196_;
  assign new_n7199_ = ~new_n7197_ & ~new_n7198_;
  assign new_n7200_ = new_n4475_ & ~new_n7199_;
  assign new_n7201_ = lo0055 & new_n5083_;
  assign new_n7202_ = ~new_n7194_ & ~new_n7200_;
  assign new_n7203_ = ~new_n7201_ & new_n7202_;
  assign new_n7204_ = new_n5070_ & ~new_n7203_;
  assign new_n7205_ = ~new_n4096_ & new_n7173_;
  assign new_n7206_ = lo0055 & ~new_n7173_;
  assign new_n7207_ = ~new_n7205_ & ~new_n7206_;
  assign new_n7208_ = new_n5090_ & ~new_n7207_;
  assign new_n7209_ = new_n3746_ & new_n7172_;
  assign new_n7210_ = ~new_n7208_ & ~new_n7209_;
  assign new_n7211_ = new_n7193_ & ~new_n7204_;
  assign new_n7212_ = new_n7210_ & new_n7211_;
  assign new_n7213_ = lo0055 & new_n5505_;
  assign new_n7214_ = lo0055 & new_n5135_;
  assign new_n7215_ = ~lo1044 & new_n7172_;
  assign new_n7216_ = new_n4007_ & new_n7215_;
  assign new_n7217_ = new_n3969_ & new_n7177_;
  assign new_n7218_ = ~new_n7216_ & ~new_n7217_;
  assign new_n7219_ = ~new_n7213_ & ~new_n7214_;
  assign new_n7220_ = new_n7218_ & new_n7219_;
  assign new_n7221_ = new_n3810_ & new_n7177_;
  assign new_n7222_ = lo0055 & new_n5112_;
  assign new_n7223_ = ~new_n7221_ & ~new_n7222_;
  assign new_n7224_ = ~new_n3879_ & new_n7223_;
  assign new_n7225_ = new_n3804_ & new_n7173_;
  assign new_n7226_ = new_n3834_ & new_n7196_;
  assign new_n7227_ = new_n3678_ & new_n7226_;
  assign new_n7228_ = new_n7224_ & ~new_n7225_;
  assign new_n7229_ = ~new_n7227_ & new_n7228_;
  assign new_n7230_ = ~new_n5105_ & new_n7177_;
  assign new_n7231_ = new_n7229_ & ~new_n7230_;
  assign new_n7232_ = new_n3815_ & new_n7172_;
  assign new_n7233_ = new_n4088_ & new_n7173_;
  assign new_n7234_ = ~new_n7232_ & ~new_n7233_;
  assign new_n7235_ = new_n3820_ & new_n7177_;
  assign new_n7236_ = new_n3870_ & new_n7215_;
  assign new_n7237_ = ~new_n7235_ & ~new_n7236_;
  assign new_n7238_ = ~new_n4069_ & new_n7173_;
  assign new_n7239_ = new_n7231_ & new_n7234_;
  assign new_n7240_ = new_n7237_ & new_n7239_;
  assign new_n7241_ = ~new_n7238_ & new_n7240_;
  assign new_n7242_ = new_n7220_ & new_n7241_;
  assign new_n7243_ = new_n4050_ & new_n7173_;
  assign new_n7244_ = lo0055 & new_n5562_;
  assign new_n7245_ = new_n3763_ & new_n7177_;
  assign new_n7246_ = new_n3780_ & new_n7173_;
  assign new_n7247_ = ~new_n7245_ & ~new_n7246_;
  assign new_n7248_ = new_n3794_ & new_n7172_;
  assign new_n7249_ = new_n7247_ & ~new_n7248_;
  assign new_n7250_ = lo0055 & new_n5155_;
  assign new_n7251_ = new_n3777_ & new_n7250_;
  assign new_n7252_ = lo0055 & ~new_n4632_;
  assign new_n7253_ = new_n5565_ & new_n7252_;
  assign new_n7254_ = ~new_n7251_ & ~new_n7253_;
  assign new_n7255_ = ~new_n5460_ & new_n7172_;
  assign new_n7256_ = new_n7254_ & ~new_n7255_;
  assign new_n7257_ = ~new_n7243_ & ~new_n7244_;
  assign new_n7258_ = new_n7249_ & new_n7257_;
  assign new_n7259_ = new_n7256_ & new_n7258_;
  assign new_n7260_ = new_n4041_ & new_n7173_;
  assign new_n7261_ = new_n7259_ & ~new_n7260_;
  assign new_n7262_ = lo0055 & ~new_n5216_;
  assign new_n7263_ = new_n4133_ & new_n7173_;
  assign new_n7264_ = ~new_n7262_ & ~new_n7263_;
  assign new_n7265_ = new_n3974_ & new_n7196_;
  assign new_n7266_ = ~new_n4135_ & new_n7265_;
  assign new_n7267_ = lo0055 & new_n5225_;
  assign new_n7268_ = new_n7264_ & ~new_n7266_;
  assign new_n7269_ = ~new_n7267_ & new_n7268_;
  assign new_n7270_ = new_n3948_ & new_n7173_;
  assign new_n7271_ = new_n7269_ & ~new_n7270_;
  assign new_n7272_ = lo0055 & ~lo0993;
  assign new_n7273_ = new_n3927_ & new_n7272_;
  assign new_n7274_ = new_n3953_ & new_n7173_;
  assign new_n7275_ = ~new_n7273_ & ~new_n7274_;
  assign new_n7276_ = lo0055 & new_n3678_;
  assign new_n7277_ = new_n3786_ & new_n7173_;
  assign new_n7278_ = new_n5139_ & new_n7276_;
  assign new_n7279_ = ~new_n7277_ & ~new_n7278_;
  assign new_n7280_ = new_n7261_ & new_n7271_;
  assign new_n7281_ = new_n7275_ & new_n7280_;
  assign new_n7282_ = new_n7279_ & new_n7281_;
  assign new_n7283_ = new_n7190_ & new_n7212_;
  assign new_n7284_ = new_n7242_ & new_n7283_;
  assign li0055 = ~new_n7282_ | ~new_n7284_;
  assign new_n7286_ = ~lo0024 & lo0056;
  assign new_n7287_ = new_n4050_ & new_n7286_;
  assign new_n7288_ = lo0056 & new_n5562_;
  assign new_n7289_ = lo0056 & ~lo0314;
  assign new_n7290_ = lo0056 & new_n5155_;
  assign new_n7291_ = new_n3777_ & new_n7290_;
  assign new_n7292_ = lo0056 & ~new_n4632_;
  assign new_n7293_ = new_n5565_ & new_n7292_;
  assign new_n7294_ = ~new_n7291_ & ~new_n7293_;
  assign new_n7295_ = ~new_n5460_ & new_n7289_;
  assign new_n7296_ = new_n7294_ & ~new_n7295_;
  assign new_n7297_ = lo0056 & ~lo0841;
  assign new_n7298_ = new_n3763_ & new_n7297_;
  assign new_n7299_ = new_n3780_ & new_n7286_;
  assign new_n7300_ = ~new_n7298_ & ~new_n7299_;
  assign new_n7301_ = new_n3794_ & new_n7289_;
  assign new_n7302_ = new_n7300_ & ~new_n7301_;
  assign new_n7303_ = ~new_n7287_ & ~new_n7288_;
  assign new_n7304_ = new_n7296_ & new_n7303_;
  assign new_n7305_ = new_n7302_ & new_n7304_;
  assign new_n7306_ = new_n4041_ & new_n7286_;
  assign new_n7307_ = new_n7305_ & ~new_n7306_;
  assign new_n7308_ = lo0056 & ~new_n5216_;
  assign new_n7309_ = ~lo0024 & ~lo0056;
  assign new_n7310_ = new_n3948_ & ~new_n7309_;
  assign new_n7311_ = lo0056 & new_n5225_;
  assign new_n7312_ = lo0056 & li0583;
  assign new_n7313_ = new_n3974_ & new_n7312_;
  assign new_n7314_ = ~new_n4135_ & new_n7313_;
  assign new_n7315_ = ~new_n7308_ & ~new_n7310_;
  assign new_n7316_ = ~new_n7311_ & new_n7315_;
  assign new_n7317_ = ~new_n7314_ & new_n7316_;
  assign new_n7318_ = new_n4133_ & new_n7286_;
  assign new_n7319_ = new_n7317_ & ~new_n7318_;
  assign new_n7320_ = lo0056 & new_n3678_;
  assign new_n7321_ = new_n3786_ & new_n7286_;
  assign new_n7322_ = new_n5139_ & new_n7320_;
  assign new_n7323_ = ~new_n7321_ & ~new_n7322_;
  assign new_n7324_ = new_n7319_ & new_n7323_;
  assign new_n7325_ = new_n7307_ & new_n7324_;
  assign new_n7326_ = new_n3804_ & new_n7286_;
  assign new_n7327_ = new_n3834_ & new_n7312_;
  assign new_n7328_ = new_n3678_ & new_n7327_;
  assign new_n7329_ = lo0056 & new_n5112_;
  assign new_n7330_ = new_n3810_ & new_n7297_;
  assign new_n7331_ = ~new_n7326_ & ~new_n7328_;
  assign new_n7332_ = ~new_n7329_ & new_n7331_;
  assign new_n7333_ = ~new_n7330_ & new_n7332_;
  assign new_n7334_ = ~new_n5105_ & new_n7297_;
  assign new_n7335_ = new_n7333_ & ~new_n7334_;
  assign new_n7336_ = new_n3815_ & new_n7289_;
  assign new_n7337_ = new_n4088_ & new_n7286_;
  assign new_n7338_ = ~new_n7336_ & ~new_n7337_;
  assign new_n7339_ = ~lo1044 & new_n7289_;
  assign new_n7340_ = new_n3820_ & new_n7297_;
  assign new_n7341_ = new_n3870_ & new_n7339_;
  assign new_n7342_ = ~new_n7340_ & ~new_n7341_;
  assign new_n7343_ = ~new_n4069_ & new_n7286_;
  assign new_n7344_ = new_n7335_ & new_n7338_;
  assign new_n7345_ = new_n7342_ & new_n7344_;
  assign new_n7346_ = ~new_n7343_ & new_n7345_;
  assign new_n7347_ = new_n7325_ & new_n7346_;
  assign new_n7348_ = lo0056 & new_n5194_;
  assign new_n7349_ = ~new_n7286_ & ~new_n7348_;
  assign new_n7350_ = new_n3936_ & ~new_n7349_;
  assign new_n7351_ = new_n3625_ & new_n7286_;
  assign new_n7352_ = ~new_n7350_ & ~new_n7351_;
  assign new_n7353_ = lo0056 & new_n3706_;
  assign new_n7354_ = lo0056 & new_n5818_;
  assign new_n7355_ = ~new_n5184_ & new_n7354_;
  assign new_n7356_ = new_n7352_ & ~new_n7353_;
  assign new_n7357_ = ~new_n7355_ & new_n7356_;
  assign new_n7358_ = ~new_n5201_ & new_n7297_;
  assign new_n7359_ = new_n7357_ & ~new_n7358_;
  assign new_n7360_ = ~new_n5060_ & new_n7289_;
  assign new_n7361_ = new_n3940_ & new_n7286_;
  assign new_n7362_ = ~new_n7360_ & ~new_n7361_;
  assign new_n7363_ = new_n7359_ & new_n7362_;
  assign new_n7364_ = new_n4020_ & new_n7286_;
  assign new_n7365_ = ~new_n5096_ & new_n7297_;
  assign new_n7366_ = ~new_n7364_ & ~new_n7365_;
  assign new_n7367_ = lo0056 & new_n5071_;
  assign new_n7368_ = lo0056 & new_n4219_;
  assign new_n7369_ = ~new_n5074_ & new_n7368_;
  assign new_n7370_ = ~new_n5076_ & new_n7312_;
  assign new_n7371_ = ~new_n7369_ & ~new_n7370_;
  assign new_n7372_ = new_n4475_ & ~new_n7371_;
  assign new_n7373_ = lo0056 & new_n5083_;
  assign new_n7374_ = ~new_n7367_ & ~new_n7372_;
  assign new_n7375_ = ~new_n7373_ & new_n7374_;
  assign new_n7376_ = new_n5070_ & ~new_n7375_;
  assign new_n7377_ = ~new_n4096_ & new_n7286_;
  assign new_n7378_ = lo0056 & ~new_n7286_;
  assign new_n7379_ = ~new_n7377_ & ~new_n7378_;
  assign new_n7380_ = new_n5090_ & ~new_n7379_;
  assign new_n7381_ = new_n3746_ & new_n7289_;
  assign new_n7382_ = ~new_n7380_ & ~new_n7381_;
  assign new_n7383_ = new_n7366_ & ~new_n7376_;
  assign new_n7384_ = new_n7382_ & new_n7383_;
  assign new_n7385_ = lo0056 & new_n5505_;
  assign new_n7386_ = lo0056 & new_n5135_;
  assign new_n7387_ = lo0056 & ~lo0993;
  assign new_n7388_ = new_n3927_ & new_n7387_;
  assign new_n7389_ = new_n3953_ & new_n7286_;
  assign new_n7390_ = ~new_n7388_ & ~new_n7389_;
  assign new_n7391_ = new_n4007_ & new_n7339_;
  assign new_n7392_ = new_n3969_ & new_n7297_;
  assign new_n7393_ = ~new_n7391_ & ~new_n7392_;
  assign new_n7394_ = ~new_n7385_ & ~new_n7386_;
  assign new_n7395_ = new_n7390_ & new_n7394_;
  assign new_n7396_ = new_n7393_ & new_n7395_;
  assign new_n7397_ = new_n7347_ & new_n7363_;
  assign new_n7398_ = new_n7384_ & new_n7397_;
  assign li0056 = ~new_n7396_ | ~new_n7398_;
  assign new_n7400_ = lo0057 & ~lo0841;
  assign new_n7401_ = ~lo0024 & lo0057;
  assign new_n7402_ = new_n4020_ & new_n7401_;
  assign new_n7403_ = ~new_n5096_ & new_n7400_;
  assign new_n7404_ = ~new_n7402_ & ~new_n7403_;
  assign new_n7405_ = lo0057 & new_n5071_;
  assign new_n7406_ = lo0057 & new_n4219_;
  assign new_n7407_ = lo0057 & li0583;
  assign new_n7408_ = ~new_n5074_ & new_n7406_;
  assign new_n7409_ = ~new_n5076_ & new_n7407_;
  assign new_n7410_ = ~new_n7408_ & ~new_n7409_;
  assign new_n7411_ = new_n4475_ & ~new_n7410_;
  assign new_n7412_ = lo0057 & new_n5083_;
  assign new_n7413_ = ~new_n7405_ & ~new_n7411_;
  assign new_n7414_ = ~new_n7412_ & new_n7413_;
  assign new_n7415_ = new_n5070_ & ~new_n7414_;
  assign new_n7416_ = ~new_n4096_ & new_n7401_;
  assign new_n7417_ = lo0057 & ~new_n7401_;
  assign new_n7418_ = ~new_n7416_ & ~new_n7417_;
  assign new_n7419_ = lo0057 & ~lo0314;
  assign new_n7420_ = new_n5090_ & ~new_n7418_;
  assign new_n7421_ = new_n3746_ & new_n7419_;
  assign new_n7422_ = ~new_n7420_ & ~new_n7421_;
  assign new_n7423_ = new_n7404_ & ~new_n7415_;
  assign new_n7424_ = new_n7422_ & new_n7423_;
  assign new_n7425_ = new_n3804_ & new_n7401_;
  assign new_n7426_ = new_n3834_ & new_n7407_;
  assign new_n7427_ = new_n3678_ & new_n7426_;
  assign new_n7428_ = lo0057 & new_n5112_;
  assign new_n7429_ = new_n3810_ & new_n7400_;
  assign new_n7430_ = ~new_n7425_ & ~new_n7427_;
  assign new_n7431_ = ~new_n7428_ & new_n7430_;
  assign new_n7432_ = ~new_n7429_ & new_n7431_;
  assign new_n7433_ = ~new_n5105_ & new_n7400_;
  assign new_n7434_ = new_n7432_ & ~new_n7433_;
  assign new_n7435_ = new_n3815_ & new_n7419_;
  assign new_n7436_ = new_n4088_ & new_n7401_;
  assign new_n7437_ = ~new_n7435_ & ~new_n7436_;
  assign new_n7438_ = ~lo1044 & new_n7419_;
  assign new_n7439_ = new_n3820_ & new_n7400_;
  assign new_n7440_ = new_n3870_ & new_n7438_;
  assign new_n7441_ = ~new_n7439_ & ~new_n7440_;
  assign new_n7442_ = ~new_n4069_ & new_n7401_;
  assign new_n7443_ = new_n7434_ & new_n7437_;
  assign new_n7444_ = new_n7441_ & new_n7443_;
  assign new_n7445_ = ~new_n7442_ & new_n7444_;
  assign new_n7446_ = new_n7424_ & new_n7445_;
  assign new_n7447_ = lo0057 & new_n5155_;
  assign new_n7448_ = new_n3777_ & new_n7447_;
  assign new_n7449_ = lo0057 & ~new_n4632_;
  assign new_n7450_ = new_n5565_ & new_n7449_;
  assign new_n7451_ = ~new_n7448_ & ~new_n7450_;
  assign new_n7452_ = new_n3780_ & new_n7401_;
  assign new_n7453_ = new_n7451_ & ~new_n7452_;
  assign new_n7454_ = new_n3794_ & new_n7419_;
  assign new_n7455_ = new_n3914_ & new_n7419_;
  assign new_n7456_ = ~new_n7454_ & ~new_n7455_;
  assign new_n7457_ = lo0841 & ~lo0924;
  assign new_n7458_ = ~new_n7400_ & ~new_n7457_;
  assign new_n7459_ = new_n3763_ & ~new_n7458_;
  assign new_n7460_ = lo0057 & lo1076;
  assign new_n7461_ = new_n4050_ & new_n7401_;
  assign new_n7462_ = new_n3773_ & new_n7460_;
  assign new_n7463_ = ~new_n7461_ & ~new_n7462_;
  assign new_n7464_ = new_n3903_ & new_n7419_;
  assign new_n7465_ = ~new_n7459_ & new_n7463_;
  assign new_n7466_ = ~new_n7464_ & new_n7465_;
  assign new_n7467_ = new_n7456_ & new_n7466_;
  assign new_n7468_ = new_n7453_ & new_n7467_;
  assign new_n7469_ = new_n4041_ & new_n7401_;
  assign new_n7470_ = new_n7468_ & ~new_n7469_;
  assign new_n7471_ = lo0057 & new_n3678_;
  assign new_n7472_ = new_n3786_ & new_n7401_;
  assign new_n7473_ = new_n5139_ & new_n7471_;
  assign new_n7474_ = ~new_n7472_ & ~new_n7473_;
  assign new_n7475_ = new_n4007_ & new_n7438_;
  assign new_n7476_ = new_n3969_ & new_n7400_;
  assign new_n7477_ = ~new_n7475_ & ~new_n7476_;
  assign new_n7478_ = lo0057 & ~new_n5216_;
  assign new_n7479_ = new_n4133_ & new_n7401_;
  assign new_n7480_ = ~new_n7478_ & ~new_n7479_;
  assign new_n7481_ = new_n3974_ & new_n7407_;
  assign new_n7482_ = ~new_n4135_ & new_n7481_;
  assign new_n7483_ = lo0057 & new_n5225_;
  assign new_n7484_ = new_n7480_ & ~new_n7482_;
  assign new_n7485_ = ~new_n7483_ & new_n7484_;
  assign new_n7486_ = new_n3948_ & new_n7401_;
  assign new_n7487_ = new_n7485_ & ~new_n7486_;
  assign new_n7488_ = new_n7470_ & new_n7474_;
  assign new_n7489_ = new_n7477_ & new_n7488_;
  assign new_n7490_ = new_n7487_ & new_n7489_;
  assign new_n7491_ = lo0057 & new_n5505_;
  assign new_n7492_ = lo0057 & ~new_n5134_;
  assign new_n7493_ = ~new_n3714_ & ~new_n3725_;
  assign new_n7494_ = new_n7400_ & ~new_n7493_;
  assign new_n7495_ = new_n3625_ & new_n7401_;
  assign new_n7496_ = ~new_n7494_ & ~new_n7495_;
  assign new_n7497_ = ~lo0057 & ~lo0841;
  assign new_n7498_ = lo0057 & new_n5194_;
  assign new_n7499_ = ~new_n7401_ & ~new_n7498_;
  assign new_n7500_ = new_n3936_ & ~new_n7499_;
  assign new_n7501_ = new_n3931_ & ~new_n7497_;
  assign new_n7502_ = ~new_n7500_ & ~new_n7501_;
  assign new_n7503_ = lo0057 & new_n5818_;
  assign new_n7504_ = ~new_n5184_ & new_n7503_;
  assign new_n7505_ = lo0057 & new_n3706_;
  assign new_n7506_ = new_n7496_ & new_n7502_;
  assign new_n7507_ = ~new_n7504_ & new_n7506_;
  assign new_n7508_ = ~new_n7505_ & new_n7507_;
  assign new_n7509_ = new_n5133_ & new_n7492_;
  assign new_n7510_ = new_n7508_ & ~new_n7509_;
  assign new_n7511_ = ~new_n7491_ & new_n7510_;
  assign new_n7512_ = new_n7490_ & new_n7511_;
  assign new_n7513_ = ~new_n5060_ & new_n7419_;
  assign new_n7514_ = new_n3940_ & new_n7401_;
  assign new_n7515_ = ~new_n7513_ & ~new_n7514_;
  assign new_n7516_ = lo0057 & ~lo0993;
  assign new_n7517_ = new_n3927_ & new_n7516_;
  assign new_n7518_ = new_n3953_ & new_n7401_;
  assign new_n7519_ = ~new_n7517_ & ~new_n7518_;
  assign new_n7520_ = new_n7515_ & new_n7519_;
  assign new_n7521_ = new_n7446_ & new_n7512_;
  assign li0057 = ~new_n7520_ | ~new_n7521_;
  assign new_n7523_ = lo0058 & ~lo0841;
  assign new_n7524_ = ~new_n5201_ & new_n7523_;
  assign new_n7525_ = ~lo0024 & lo0058;
  assign new_n7526_ = lo0058 & new_n5194_;
  assign new_n7527_ = ~new_n7525_ & ~new_n7526_;
  assign new_n7528_ = new_n3936_ & ~new_n7527_;
  assign new_n7529_ = new_n3625_ & new_n7525_;
  assign new_n7530_ = ~new_n7528_ & ~new_n7529_;
  assign new_n7531_ = lo0058 & new_n5608_;
  assign new_n7532_ = ~new_n5184_ & new_n7531_;
  assign new_n7533_ = lo0058 & new_n3706_;
  assign new_n7534_ = ~new_n7524_ & new_n7530_;
  assign new_n7535_ = ~new_n7532_ & new_n7534_;
  assign new_n7536_ = ~new_n7533_ & new_n7535_;
  assign new_n7537_ = new_n4050_ & new_n7525_;
  assign new_n7538_ = lo0058 & new_n5562_;
  assign new_n7539_ = lo0058 & ~lo0314;
  assign new_n7540_ = lo0058 & new_n5155_;
  assign new_n7541_ = new_n3777_ & new_n7540_;
  assign new_n7542_ = lo0058 & ~new_n4632_;
  assign new_n7543_ = new_n5565_ & new_n7542_;
  assign new_n7544_ = ~new_n7541_ & ~new_n7543_;
  assign new_n7545_ = ~new_n5460_ & new_n7539_;
  assign new_n7546_ = new_n7544_ & ~new_n7545_;
  assign new_n7547_ = new_n3763_ & new_n7523_;
  assign new_n7548_ = new_n3780_ & new_n7525_;
  assign new_n7549_ = ~new_n7547_ & ~new_n7548_;
  assign new_n7550_ = new_n3794_ & new_n7539_;
  assign new_n7551_ = new_n7549_ & ~new_n7550_;
  assign new_n7552_ = ~new_n7537_ & ~new_n7538_;
  assign new_n7553_ = new_n7546_ & new_n7552_;
  assign new_n7554_ = new_n7551_ & new_n7553_;
  assign new_n7555_ = new_n4041_ & new_n7525_;
  assign new_n7556_ = new_n7554_ & ~new_n7555_;
  assign new_n7557_ = new_n7536_ & new_n7556_;
  assign new_n7558_ = lo0058 & new_n5505_;
  assign new_n7559_ = ~lo1044 & new_n7539_;
  assign new_n7560_ = new_n4007_ & new_n7559_;
  assign new_n7561_ = new_n3969_ & new_n7523_;
  assign new_n7562_ = ~new_n7560_ & ~new_n7561_;
  assign new_n7563_ = new_n3786_ & new_n7525_;
  assign new_n7564_ = lo0058 & new_n5140_;
  assign new_n7565_ = new_n3948_ & new_n7525_;
  assign new_n7566_ = ~new_n7564_ & ~new_n7565_;
  assign new_n7567_ = new_n7562_ & ~new_n7563_;
  assign new_n7568_ = new_n7566_ & new_n7567_;
  assign new_n7569_ = ~new_n4637_ & new_n7568_;
  assign new_n7570_ = new_n3804_ & new_n7525_;
  assign new_n7571_ = lo0058 & li0583;
  assign new_n7572_ = new_n3834_ & new_n7571_;
  assign new_n7573_ = new_n3678_ & new_n7572_;
  assign new_n7574_ = lo0058 & new_n5112_;
  assign new_n7575_ = new_n3810_ & new_n7523_;
  assign new_n7576_ = ~new_n7570_ & ~new_n7573_;
  assign new_n7577_ = ~new_n7574_ & new_n7576_;
  assign new_n7578_ = ~new_n7575_ & new_n7577_;
  assign new_n7579_ = new_n3815_ & new_n7539_;
  assign new_n7580_ = new_n7578_ & ~new_n7579_;
  assign new_n7581_ = ~new_n4069_ & new_n7525_;
  assign new_n7582_ = new_n3820_ & new_n7523_;
  assign new_n7583_ = new_n3870_ & new_n7559_;
  assign new_n7584_ = ~new_n7582_ & ~new_n7583_;
  assign new_n7585_ = new_n7580_ & ~new_n7581_;
  assign new_n7586_ = new_n7584_ & new_n7585_;
  assign new_n7587_ = lo0058 & new_n3857_;
  assign new_n7588_ = new_n7586_ & ~new_n7587_;
  assign new_n7589_ = ~new_n5104_ & new_n7523_;
  assign new_n7590_ = new_n4088_ & new_n7525_;
  assign new_n7591_ = ~new_n7589_ & ~new_n7590_;
  assign new_n7592_ = new_n7588_ & new_n7591_;
  assign new_n7593_ = new_n7569_ & new_n7592_;
  assign new_n7594_ = lo0058 & ~new_n5134_;
  assign new_n7595_ = new_n3974_ & new_n7571_;
  assign new_n7596_ = ~new_n4135_ & new_n7595_;
  assign new_n7597_ = lo0058 & new_n5225_;
  assign new_n7598_ = ~new_n7596_ & ~new_n7597_;
  assign new_n7599_ = lo0058 & ~new_n5216_;
  assign new_n7600_ = new_n4133_ & new_n7525_;
  assign new_n7601_ = ~new_n7599_ & ~new_n7600_;
  assign new_n7602_ = new_n7598_ & new_n7601_;
  assign new_n7603_ = new_n5133_ & new_n7594_;
  assign new_n7604_ = new_n7602_ & ~new_n7603_;
  assign new_n7605_ = new_n7557_ & ~new_n7558_;
  assign new_n7606_ = new_n7593_ & new_n7605_;
  assign new_n7607_ = new_n7604_ & new_n7606_;
  assign new_n7608_ = ~new_n5060_ & new_n7539_;
  assign new_n7609_ = new_n3940_ & new_n7525_;
  assign new_n7610_ = ~new_n7608_ & ~new_n7609_;
  assign new_n7611_ = lo0058 & ~lo0993;
  assign new_n7612_ = new_n3927_ & new_n7611_;
  assign new_n7613_ = new_n3953_ & new_n7525_;
  assign new_n7614_ = ~new_n7612_ & ~new_n7613_;
  assign new_n7615_ = lo0058 & new_n5071_;
  assign new_n7616_ = lo0058 & new_n4219_;
  assign new_n7617_ = ~new_n5074_ & new_n7616_;
  assign new_n7618_ = ~new_n5076_ & new_n7571_;
  assign new_n7619_ = ~new_n7617_ & ~new_n7618_;
  assign new_n7620_ = new_n4475_ & ~new_n7619_;
  assign new_n7621_ = lo0058 & new_n5083_;
  assign new_n7622_ = ~new_n7615_ & ~new_n7620_;
  assign new_n7623_ = ~new_n7621_ & new_n7622_;
  assign new_n7624_ = new_n3746_ & new_n7539_;
  assign new_n7625_ = ~new_n4096_ & new_n7525_;
  assign new_n7626_ = lo0058 & ~new_n7525_;
  assign new_n7627_ = ~new_n7625_ & ~new_n7626_;
  assign new_n7628_ = new_n5090_ & ~new_n7627_;
  assign new_n7629_ = ~new_n7624_ & ~new_n7628_;
  assign new_n7630_ = new_n5070_ & ~new_n7623_;
  assign new_n7631_ = new_n7629_ & ~new_n7630_;
  assign new_n7632_ = new_n4020_ & new_n7525_;
  assign new_n7633_ = ~new_n5096_ & new_n7523_;
  assign new_n7634_ = ~new_n7632_ & ~new_n7633_;
  assign new_n7635_ = new_n7610_ & new_n7614_;
  assign new_n7636_ = new_n7631_ & new_n7635_;
  assign new_n7637_ = new_n7634_ & new_n7636_;
  assign li0058 = ~new_n7607_ | ~new_n7637_;
  assign new_n7639_ = lo0059 & new_n5135_;
  assign new_n7640_ = lo0059 & ~lo0841;
  assign new_n7641_ = lo0059 & ~lo0314;
  assign new_n7642_ = ~lo1044 & new_n7641_;
  assign new_n7643_ = new_n4007_ & new_n7642_;
  assign new_n7644_ = new_n3969_ & new_n7640_;
  assign new_n7645_ = ~new_n7643_ & ~new_n7644_;
  assign new_n7646_ = ~new_n7639_ & new_n7645_;
  assign new_n7647_ = lo0059 & new_n5505_;
  assign new_n7648_ = lo0059 & ~lo0993;
  assign new_n7649_ = ~lo0024 & lo0059;
  assign new_n7650_ = new_n3927_ & new_n7648_;
  assign new_n7651_ = new_n3953_ & new_n7649_;
  assign new_n7652_ = ~new_n7650_ & ~new_n7651_;
  assign new_n7653_ = new_n7646_ & ~new_n7647_;
  assign new_n7654_ = new_n7652_ & new_n7653_;
  assign new_n7655_ = new_n4020_ & new_n7649_;
  assign new_n7656_ = ~new_n5096_ & new_n7640_;
  assign new_n7657_ = ~new_n7655_ & ~new_n7656_;
  assign new_n7658_ = lo0059 & new_n5071_;
  assign new_n7659_ = lo0059 & new_n4219_;
  assign new_n7660_ = lo0059 & li0583;
  assign new_n7661_ = ~new_n5074_ & new_n7659_;
  assign new_n7662_ = ~new_n5076_ & new_n7660_;
  assign new_n7663_ = ~new_n7661_ & ~new_n7662_;
  assign new_n7664_ = new_n4475_ & ~new_n7663_;
  assign new_n7665_ = lo0059 & new_n5083_;
  assign new_n7666_ = ~new_n7658_ & ~new_n7664_;
  assign new_n7667_ = ~new_n7665_ & new_n7666_;
  assign new_n7668_ = new_n5070_ & ~new_n7667_;
  assign new_n7669_ = ~new_n4096_ & new_n7649_;
  assign new_n7670_ = lo0059 & ~new_n7649_;
  assign new_n7671_ = ~new_n7669_ & ~new_n7670_;
  assign new_n7672_ = new_n5090_ & ~new_n7671_;
  assign new_n7673_ = new_n3746_ & new_n7641_;
  assign new_n7674_ = ~new_n7672_ & ~new_n7673_;
  assign new_n7675_ = new_n7657_ & ~new_n7668_;
  assign new_n7676_ = new_n7674_ & new_n7675_;
  assign new_n7677_ = new_n7654_ & new_n7676_;
  assign new_n7678_ = ~new_n5060_ & new_n7641_;
  assign new_n7679_ = new_n3940_ & new_n7649_;
  assign new_n7680_ = ~new_n7678_ & ~new_n7679_;
  assign new_n7681_ = lo0059 & new_n5194_;
  assign new_n7682_ = ~new_n7649_ & ~new_n7681_;
  assign new_n7683_ = new_n3936_ & ~new_n7682_;
  assign new_n7684_ = new_n3625_ & new_n7649_;
  assign new_n7685_ = ~new_n7683_ & ~new_n7684_;
  assign new_n7686_ = lo0059 & new_n3706_;
  assign new_n7687_ = lo0059 & new_n5818_;
  assign new_n7688_ = ~new_n5184_ & new_n7687_;
  assign new_n7689_ = new_n7685_ & ~new_n7686_;
  assign new_n7690_ = ~new_n7688_ & new_n7689_;
  assign new_n7691_ = ~new_n5201_ & new_n7640_;
  assign new_n7692_ = new_n7690_ & ~new_n7691_;
  assign new_n7693_ = new_n7680_ & new_n7692_;
  assign new_n7694_ = lo0059 & lo1076;
  assign new_n7695_ = new_n3773_ & new_n7694_;
  assign new_n7696_ = new_n4050_ & new_n7649_;
  assign new_n7697_ = ~new_n7695_ & ~new_n7696_;
  assign new_n7698_ = new_n3794_ & new_n7641_;
  assign new_n7699_ = new_n3780_ & new_n7649_;
  assign new_n7700_ = ~new_n7698_ & ~new_n7699_;
  assign new_n7701_ = new_n3914_ & new_n7641_;
  assign new_n7702_ = new_n7700_ & ~new_n7701_;
  assign new_n7703_ = lo0841 & lo0924;
  assign new_n7704_ = ~new_n7640_ & ~new_n7703_;
  assign new_n7705_ = new_n3763_ & ~new_n7704_;
  assign new_n7706_ = lo0059 & new_n5155_;
  assign new_n7707_ = new_n3777_ & new_n7706_;
  assign new_n7708_ = lo0059 & ~new_n4632_;
  assign new_n7709_ = new_n5565_ & new_n7708_;
  assign new_n7710_ = ~new_n7707_ & ~new_n7709_;
  assign new_n7711_ = new_n3903_ & new_n7641_;
  assign new_n7712_ = new_n7710_ & ~new_n7711_;
  assign new_n7713_ = new_n7697_ & new_n7702_;
  assign new_n7714_ = ~new_n7705_ & new_n7713_;
  assign new_n7715_ = new_n7712_ & new_n7714_;
  assign new_n7716_ = new_n4041_ & new_n7649_;
  assign new_n7717_ = new_n7715_ & ~new_n7716_;
  assign new_n7718_ = lo0059 & ~new_n5216_;
  assign new_n7719_ = new_n4133_ & new_n7649_;
  assign new_n7720_ = ~new_n7718_ & ~new_n7719_;
  assign new_n7721_ = new_n3974_ & new_n7660_;
  assign new_n7722_ = ~new_n4135_ & new_n7721_;
  assign new_n7723_ = lo0059 & new_n5225_;
  assign new_n7724_ = new_n7720_ & ~new_n7722_;
  assign new_n7725_ = ~new_n7723_ & new_n7724_;
  assign new_n7726_ = new_n3948_ & new_n7649_;
  assign new_n7727_ = new_n7725_ & ~new_n7726_;
  assign new_n7728_ = lo0059 & new_n3678_;
  assign new_n7729_ = new_n3786_ & new_n7649_;
  assign new_n7730_ = new_n5139_ & new_n7728_;
  assign new_n7731_ = ~new_n7729_ & ~new_n7730_;
  assign new_n7732_ = new_n7727_ & new_n7731_;
  assign new_n7733_ = new_n7717_ & new_n7732_;
  assign new_n7734_ = new_n3804_ & new_n7649_;
  assign new_n7735_ = new_n3834_ & new_n7660_;
  assign new_n7736_ = new_n3678_ & new_n7735_;
  assign new_n7737_ = lo0059 & new_n5112_;
  assign new_n7738_ = new_n3810_ & new_n7640_;
  assign new_n7739_ = ~new_n7734_ & ~new_n7736_;
  assign new_n7740_ = ~new_n7737_ & new_n7739_;
  assign new_n7741_ = ~new_n7738_ & new_n7740_;
  assign new_n7742_ = ~new_n5105_ & new_n7640_;
  assign new_n7743_ = new_n7741_ & ~new_n7742_;
  assign new_n7744_ = new_n3815_ & new_n7641_;
  assign new_n7745_ = new_n4088_ & new_n7649_;
  assign new_n7746_ = ~new_n7744_ & ~new_n7745_;
  assign new_n7747_ = new_n3820_ & new_n7640_;
  assign new_n7748_ = new_n3870_ & new_n7642_;
  assign new_n7749_ = ~new_n7747_ & ~new_n7748_;
  assign new_n7750_ = ~new_n4069_ & new_n7649_;
  assign new_n7751_ = new_n7743_ & new_n7746_;
  assign new_n7752_ = new_n7749_ & new_n7751_;
  assign new_n7753_ = ~new_n7750_ & new_n7752_;
  assign new_n7754_ = new_n7733_ & new_n7753_;
  assign new_n7755_ = new_n7677_ & new_n7693_;
  assign li0059 = ~new_n7754_ | ~new_n7755_;
  assign new_n7757_ = lo0060 & new_n5135_;
  assign new_n7758_ = lo0060 & ~lo0841;
  assign new_n7759_ = lo0060 & ~lo0314;
  assign new_n7760_ = ~lo1044 & new_n7759_;
  assign new_n7761_ = new_n4007_ & new_n7760_;
  assign new_n7762_ = new_n3969_ & new_n7758_;
  assign new_n7763_ = ~new_n7761_ & ~new_n7762_;
  assign new_n7764_ = ~new_n7757_ & new_n7763_;
  assign new_n7765_ = lo0060 & new_n5505_;
  assign new_n7766_ = lo0060 & ~lo0993;
  assign new_n7767_ = ~lo0024 & lo0060;
  assign new_n7768_ = new_n3927_ & new_n7766_;
  assign new_n7769_ = new_n3953_ & new_n7767_;
  assign new_n7770_ = ~new_n7768_ & ~new_n7769_;
  assign new_n7771_ = new_n7764_ & ~new_n7765_;
  assign new_n7772_ = new_n7770_ & new_n7771_;
  assign new_n7773_ = new_n4020_ & new_n7767_;
  assign new_n7774_ = ~new_n5096_ & new_n7758_;
  assign new_n7775_ = ~new_n7773_ & ~new_n7774_;
  assign new_n7776_ = ~new_n4096_ & new_n7767_;
  assign new_n7777_ = lo0060 & ~new_n7767_;
  assign new_n7778_ = ~new_n7776_ & ~new_n7777_;
  assign new_n7779_ = new_n5090_ & ~new_n7778_;
  assign new_n7780_ = new_n3746_ & new_n7759_;
  assign new_n7781_ = ~new_n7779_ & ~new_n7780_;
  assign new_n7782_ = ~new_n4421_ & ~new_n6950_;
  assign new_n7783_ = lo0060 & li0583;
  assign new_n7784_ = ~new_n5076_ & new_n7783_;
  assign new_n7785_ = lo0060 & new_n5545_;
  assign new_n7786_ = ~new_n4421_ & new_n4475_;
  assign new_n7787_ = ~new_n7784_ & ~new_n7785_;
  assign new_n7788_ = new_n7786_ & ~new_n7787_;
  assign new_n7789_ = lo0060 & new_n7782_;
  assign new_n7790_ = ~new_n7788_ & ~new_n7789_;
  assign new_n7791_ = ~new_n4421_ & new_n4423_;
  assign new_n7792_ = new_n7790_ & ~new_n7791_;
  assign new_n7793_ = new_n3612_ & ~new_n7792_;
  assign new_n7794_ = new_n4524_ & new_n7793_;
  assign new_n7795_ = new_n7775_ & new_n7781_;
  assign new_n7796_ = ~new_n7794_ & new_n7795_;
  assign new_n7797_ = new_n7772_ & new_n7796_;
  assign new_n7798_ = ~new_n5060_ & new_n7759_;
  assign new_n7799_ = new_n3940_ & new_n7767_;
  assign new_n7800_ = ~new_n7798_ & ~new_n7799_;
  assign new_n7801_ = lo0060 & new_n5194_;
  assign new_n7802_ = ~new_n7767_ & ~new_n7801_;
  assign new_n7803_ = new_n3936_ & ~new_n7802_;
  assign new_n7804_ = new_n3625_ & new_n7767_;
  assign new_n7805_ = ~new_n7803_ & ~new_n7804_;
  assign new_n7806_ = lo0060 & new_n3706_;
  assign new_n7807_ = lo0060 & new_n5818_;
  assign new_n7808_ = ~new_n5184_ & new_n7807_;
  assign new_n7809_ = new_n7805_ & ~new_n7806_;
  assign new_n7810_ = ~new_n7808_ & new_n7809_;
  assign new_n7811_ = ~new_n5201_ & new_n7758_;
  assign new_n7812_ = new_n7810_ & ~new_n7811_;
  assign new_n7813_ = new_n7800_ & new_n7812_;
  assign new_n7814_ = new_n4050_ & new_n7767_;
  assign new_n7815_ = lo0060 & new_n5562_;
  assign new_n7816_ = lo0060 & new_n5155_;
  assign new_n7817_ = new_n3777_ & new_n7816_;
  assign new_n7818_ = lo0060 & ~new_n4632_;
  assign new_n7819_ = new_n5565_ & new_n7818_;
  assign new_n7820_ = ~new_n7817_ & ~new_n7819_;
  assign new_n7821_ = ~new_n5460_ & new_n7759_;
  assign new_n7822_ = new_n7820_ & ~new_n7821_;
  assign new_n7823_ = new_n3763_ & new_n7758_;
  assign new_n7824_ = new_n3780_ & new_n7767_;
  assign new_n7825_ = ~new_n7823_ & ~new_n7824_;
  assign new_n7826_ = new_n3794_ & new_n7759_;
  assign new_n7827_ = new_n7825_ & ~new_n7826_;
  assign new_n7828_ = ~new_n7814_ & ~new_n7815_;
  assign new_n7829_ = new_n7822_ & new_n7828_;
  assign new_n7830_ = new_n7827_ & new_n7829_;
  assign new_n7831_ = new_n4041_ & new_n7767_;
  assign new_n7832_ = new_n7830_ & ~new_n7831_;
  assign new_n7833_ = lo0060 & ~new_n5216_;
  assign new_n7834_ = new_n4133_ & new_n7767_;
  assign new_n7835_ = ~new_n7833_ & ~new_n7834_;
  assign new_n7836_ = new_n3974_ & new_n7783_;
  assign new_n7837_ = ~new_n4135_ & new_n7836_;
  assign new_n7838_ = lo0060 & new_n5225_;
  assign new_n7839_ = new_n7835_ & ~new_n7837_;
  assign new_n7840_ = ~new_n7838_ & new_n7839_;
  assign new_n7841_ = new_n3948_ & new_n7767_;
  assign new_n7842_ = new_n7840_ & ~new_n7841_;
  assign new_n7843_ = lo0060 & new_n3678_;
  assign new_n7844_ = new_n3786_ & new_n7767_;
  assign new_n7845_ = new_n5139_ & new_n7843_;
  assign new_n7846_ = ~new_n7844_ & ~new_n7845_;
  assign new_n7847_ = new_n7842_ & new_n7846_;
  assign new_n7848_ = new_n7832_ & new_n7847_;
  assign new_n7849_ = new_n3804_ & new_n7767_;
  assign new_n7850_ = new_n3834_ & new_n7783_;
  assign new_n7851_ = new_n3678_ & new_n7850_;
  assign new_n7852_ = lo0060 & new_n5112_;
  assign new_n7853_ = new_n3810_ & new_n7758_;
  assign new_n7854_ = ~new_n7849_ & ~new_n7851_;
  assign new_n7855_ = ~new_n7852_ & new_n7854_;
  assign new_n7856_ = ~new_n7853_ & new_n7855_;
  assign new_n7857_ = ~new_n5105_ & new_n7758_;
  assign new_n7858_ = new_n7856_ & ~new_n7857_;
  assign new_n7859_ = new_n3815_ & new_n7759_;
  assign new_n7860_ = new_n4088_ & new_n7767_;
  assign new_n7861_ = ~new_n7859_ & ~new_n7860_;
  assign new_n7862_ = new_n3820_ & new_n7758_;
  assign new_n7863_ = new_n3870_ & new_n7760_;
  assign new_n7864_ = ~new_n7862_ & ~new_n7863_;
  assign new_n7865_ = ~new_n4069_ & new_n7767_;
  assign new_n7866_ = new_n7858_ & new_n7861_;
  assign new_n7867_ = new_n7864_ & new_n7866_;
  assign new_n7868_ = ~new_n7865_ & new_n7867_;
  assign new_n7869_ = new_n7848_ & new_n7868_;
  assign new_n7870_ = new_n7797_ & new_n7813_;
  assign li0060 = ~new_n7869_ | ~new_n7870_;
  assign new_n7872_ = lo0061 & ~lo0314;
  assign new_n7873_ = ~lo0024 & lo0061;
  assign new_n7874_ = ~new_n5060_ & new_n7872_;
  assign new_n7875_ = new_n3940_ & new_n7873_;
  assign new_n7876_ = ~new_n7874_ & ~new_n7875_;
  assign new_n7877_ = lo0061 & ~lo0841;
  assign new_n7878_ = lo0061 & new_n5194_;
  assign new_n7879_ = ~new_n7873_ & ~new_n7878_;
  assign new_n7880_ = new_n3936_ & ~new_n7879_;
  assign new_n7881_ = new_n3625_ & new_n7873_;
  assign new_n7882_ = ~new_n7880_ & ~new_n7881_;
  assign new_n7883_ = lo0061 & new_n3706_;
  assign new_n7884_ = lo0061 & new_n5818_;
  assign new_n7885_ = ~new_n5184_ & new_n7884_;
  assign new_n7886_ = new_n7882_ & ~new_n7883_;
  assign new_n7887_ = ~new_n7885_ & new_n7886_;
  assign new_n7888_ = ~new_n5201_ & new_n7877_;
  assign new_n7889_ = new_n7887_ & ~new_n7888_;
  assign new_n7890_ = new_n7876_ & new_n7889_;
  assign new_n7891_ = new_n4020_ & new_n7873_;
  assign new_n7892_ = ~new_n5096_ & new_n7877_;
  assign new_n7893_ = ~new_n7891_ & ~new_n7892_;
  assign new_n7894_ = lo0061 & new_n5071_;
  assign new_n7895_ = lo0061 & new_n4219_;
  assign new_n7896_ = lo0061 & li0583;
  assign new_n7897_ = ~new_n5074_ & new_n7895_;
  assign new_n7898_ = ~new_n5076_ & new_n7896_;
  assign new_n7899_ = ~new_n7897_ & ~new_n7898_;
  assign new_n7900_ = new_n4475_ & ~new_n7899_;
  assign new_n7901_ = lo0061 & new_n5083_;
  assign new_n7902_ = ~new_n7894_ & ~new_n7900_;
  assign new_n7903_ = ~new_n7901_ & new_n7902_;
  assign new_n7904_ = new_n5070_ & ~new_n7903_;
  assign new_n7905_ = ~new_n4096_ & new_n7873_;
  assign new_n7906_ = lo0061 & ~new_n7873_;
  assign new_n7907_ = ~new_n7905_ & ~new_n7906_;
  assign new_n7908_ = new_n5090_ & ~new_n7907_;
  assign new_n7909_ = new_n3746_ & new_n7872_;
  assign new_n7910_ = ~new_n7908_ & ~new_n7909_;
  assign new_n7911_ = new_n7893_ & ~new_n7904_;
  assign new_n7912_ = new_n7910_ & new_n7911_;
  assign new_n7913_ = lo0061 & new_n5505_;
  assign new_n7914_ = lo0061 & new_n5135_;
  assign new_n7915_ = ~lo1044 & new_n7872_;
  assign new_n7916_ = new_n4007_ & new_n7915_;
  assign new_n7917_ = new_n3969_ & new_n7877_;
  assign new_n7918_ = ~new_n7916_ & ~new_n7917_;
  assign new_n7919_ = ~new_n7913_ & ~new_n7914_;
  assign new_n7920_ = new_n7918_ & new_n7919_;
  assign new_n7921_ = new_n3804_ & new_n7873_;
  assign new_n7922_ = new_n3834_ & new_n7896_;
  assign new_n7923_ = new_n3678_ & new_n7922_;
  assign new_n7924_ = lo0061 & new_n5112_;
  assign new_n7925_ = new_n3810_ & new_n7877_;
  assign new_n7926_ = ~new_n7921_ & ~new_n7923_;
  assign new_n7927_ = ~new_n7924_ & new_n7926_;
  assign new_n7928_ = ~new_n7925_ & new_n7927_;
  assign new_n7929_ = ~new_n5105_ & new_n7877_;
  assign new_n7930_ = new_n7928_ & ~new_n7929_;
  assign new_n7931_ = new_n3815_ & new_n7872_;
  assign new_n7932_ = new_n4088_ & new_n7873_;
  assign new_n7933_ = ~new_n7931_ & ~new_n7932_;
  assign new_n7934_ = new_n3820_ & new_n7877_;
  assign new_n7935_ = new_n3870_ & new_n7915_;
  assign new_n7936_ = ~new_n7934_ & ~new_n7935_;
  assign new_n7937_ = ~new_n4069_ & new_n7873_;
  assign new_n7938_ = new_n7930_ & new_n7933_;
  assign new_n7939_ = new_n7936_ & new_n7938_;
  assign new_n7940_ = ~new_n7937_ & new_n7939_;
  assign new_n7941_ = new_n7920_ & new_n7940_;
  assign new_n7942_ = ~lo0024 & ~lo0061;
  assign new_n7943_ = new_n3786_ & ~new_n7942_;
  assign new_n7944_ = lo0061 & new_n5562_;
  assign new_n7945_ = lo0061 & new_n5155_;
  assign new_n7946_ = new_n3777_ & new_n7945_;
  assign new_n7947_ = lo0061 & ~new_n4632_;
  assign new_n7948_ = new_n5565_ & new_n7947_;
  assign new_n7949_ = ~new_n7946_ & ~new_n7948_;
  assign new_n7950_ = ~new_n5460_ & new_n7872_;
  assign new_n7951_ = new_n7949_ & ~new_n7950_;
  assign new_n7952_ = new_n3780_ & new_n7873_;
  assign new_n7953_ = new_n3763_ & new_n7877_;
  assign new_n7954_ = ~new_n7952_ & ~new_n7953_;
  assign new_n7955_ = new_n3794_ & new_n7872_;
  assign new_n7956_ = ~new_n7944_ & new_n7951_;
  assign new_n7957_ = new_n7954_ & new_n7956_;
  assign new_n7958_ = ~new_n7955_ & new_n7957_;
  assign new_n7959_ = ~new_n7943_ & new_n7958_;
  assign new_n7960_ = lo0061 & ~new_n5216_;
  assign new_n7961_ = new_n4133_ & new_n7873_;
  assign new_n7962_ = ~new_n7960_ & ~new_n7961_;
  assign new_n7963_ = new_n3974_ & new_n7896_;
  assign new_n7964_ = ~new_n4135_ & new_n7963_;
  assign new_n7965_ = lo0061 & new_n5225_;
  assign new_n7966_ = new_n7962_ & ~new_n7964_;
  assign new_n7967_ = ~new_n7965_ & new_n7966_;
  assign new_n7968_ = new_n3948_ & new_n7873_;
  assign new_n7969_ = new_n7967_ & ~new_n7968_;
  assign new_n7970_ = lo0061 & new_n5140_;
  assign new_n7971_ = new_n4041_ & new_n7873_;
  assign new_n7972_ = ~new_n7970_ & ~new_n7971_;
  assign new_n7973_ = new_n4050_ & new_n7873_;
  assign new_n7974_ = new_n7972_ & ~new_n7973_;
  assign new_n7975_ = lo0061 & ~lo0993;
  assign new_n7976_ = new_n3927_ & new_n7975_;
  assign new_n7977_ = new_n3953_ & new_n7873_;
  assign new_n7978_ = ~new_n7976_ & ~new_n7977_;
  assign new_n7979_ = new_n7959_ & new_n7969_;
  assign new_n7980_ = new_n7974_ & new_n7979_;
  assign new_n7981_ = new_n7978_ & new_n7980_;
  assign new_n7982_ = new_n7890_ & new_n7912_;
  assign new_n7983_ = new_n7941_ & new_n7982_;
  assign li0061 = ~new_n7981_ | ~new_n7983_;
  assign new_n7985_ = lo0062 & ~lo0314;
  assign new_n7986_ = ~lo0024 & lo0062;
  assign new_n7987_ = ~new_n5060_ & new_n7985_;
  assign new_n7988_ = new_n3940_ & new_n7986_;
  assign new_n7989_ = ~new_n7987_ & ~new_n7988_;
  assign new_n7990_ = lo0062 & ~lo0841;
  assign new_n7991_ = lo0062 & new_n5194_;
  assign new_n7992_ = ~new_n7986_ & ~new_n7991_;
  assign new_n7993_ = new_n3936_ & ~new_n7992_;
  assign new_n7994_ = new_n3625_ & new_n7986_;
  assign new_n7995_ = ~new_n7993_ & ~new_n7994_;
  assign new_n7996_ = lo0062 & new_n3706_;
  assign new_n7997_ = lo0062 & new_n5818_;
  assign new_n7998_ = ~new_n5184_ & new_n7997_;
  assign new_n7999_ = new_n7995_ & ~new_n7996_;
  assign new_n8000_ = ~new_n7998_ & new_n7999_;
  assign new_n8001_ = ~new_n5201_ & new_n7990_;
  assign new_n8002_ = new_n8000_ & ~new_n8001_;
  assign new_n8003_ = new_n7989_ & new_n8002_;
  assign new_n8004_ = new_n4020_ & new_n7986_;
  assign new_n8005_ = ~new_n5096_ & new_n7990_;
  assign new_n8006_ = ~new_n8004_ & ~new_n8005_;
  assign new_n8007_ = lo0062 & new_n5071_;
  assign new_n8008_ = lo0062 & new_n4219_;
  assign new_n8009_ = lo0062 & li0583;
  assign new_n8010_ = ~new_n5074_ & new_n8008_;
  assign new_n8011_ = ~new_n5076_ & new_n8009_;
  assign new_n8012_ = ~new_n8010_ & ~new_n8011_;
  assign new_n8013_ = new_n4475_ & ~new_n8012_;
  assign new_n8014_ = lo0062 & new_n5083_;
  assign new_n8015_ = ~new_n8007_ & ~new_n8013_;
  assign new_n8016_ = ~new_n8014_ & new_n8015_;
  assign new_n8017_ = new_n5070_ & ~new_n8016_;
  assign new_n8018_ = ~new_n4096_ & new_n7986_;
  assign new_n8019_ = lo0062 & ~new_n7986_;
  assign new_n8020_ = ~new_n8018_ & ~new_n8019_;
  assign new_n8021_ = new_n5090_ & ~new_n8020_;
  assign new_n8022_ = new_n3746_ & new_n7985_;
  assign new_n8023_ = ~new_n8021_ & ~new_n8022_;
  assign new_n8024_ = new_n8006_ & ~new_n8017_;
  assign new_n8025_ = new_n8023_ & new_n8024_;
  assign new_n8026_ = lo0062 & ~new_n5216_;
  assign new_n8027_ = new_n4133_ & new_n7986_;
  assign new_n8028_ = ~new_n8026_ & ~new_n8027_;
  assign new_n8029_ = new_n3974_ & new_n8009_;
  assign new_n8030_ = ~new_n4135_ & new_n8029_;
  assign new_n8031_ = lo0062 & new_n5225_;
  assign new_n8032_ = new_n8028_ & ~new_n8030_;
  assign new_n8033_ = ~new_n8031_ & new_n8032_;
  assign new_n8034_ = new_n3948_ & new_n7986_;
  assign new_n8035_ = new_n8033_ & ~new_n8034_;
  assign new_n8036_ = ~lo1044 & new_n7985_;
  assign new_n8037_ = new_n4007_ & new_n8036_;
  assign new_n8038_ = new_n3969_ & new_n7990_;
  assign new_n8039_ = ~new_n8037_ & ~new_n8038_;
  assign new_n8040_ = new_n8035_ & new_n8039_;
  assign new_n8041_ = lo0062 & new_n5562_;
  assign new_n8042_ = lo0062 & new_n5155_;
  assign new_n8043_ = new_n3777_ & new_n8042_;
  assign new_n8044_ = lo0062 & ~new_n4632_;
  assign new_n8045_ = new_n5565_ & new_n8044_;
  assign new_n8046_ = ~new_n8043_ & ~new_n8045_;
  assign new_n8047_ = ~new_n5460_ & new_n7985_;
  assign new_n8048_ = new_n8046_ & ~new_n8047_;
  assign new_n8049_ = new_n3780_ & new_n7986_;
  assign new_n8050_ = new_n3763_ & new_n7990_;
  assign new_n8051_ = ~new_n8049_ & ~new_n8050_;
  assign new_n8052_ = new_n3794_ & new_n7985_;
  assign new_n8053_ = ~new_n8041_ & new_n8048_;
  assign new_n8054_ = new_n8051_ & new_n8053_;
  assign new_n8055_ = ~new_n8052_ & new_n8054_;
  assign new_n8056_ = lo0062 & new_n4041_;
  assign new_n8057_ = new_n8055_ & ~new_n8056_;
  assign new_n8058_ = lo0062 & new_n5140_;
  assign new_n8059_ = new_n3786_ & new_n7986_;
  assign new_n8060_ = ~new_n8058_ & ~new_n8059_;
  assign new_n8061_ = new_n4050_ & new_n7986_;
  assign new_n8062_ = new_n8060_ & ~new_n8061_;
  assign new_n8063_ = new_n8040_ & new_n8057_;
  assign new_n8064_ = new_n8062_ & new_n8063_;
  assign new_n8065_ = new_n3804_ & new_n7986_;
  assign new_n8066_ = new_n3834_ & new_n8009_;
  assign new_n8067_ = new_n3678_ & new_n8066_;
  assign new_n8068_ = lo0062 & new_n5112_;
  assign new_n8069_ = new_n3810_ & new_n7990_;
  assign new_n8070_ = ~new_n8065_ & ~new_n8067_;
  assign new_n8071_ = ~new_n8068_ & new_n8070_;
  assign new_n8072_ = ~new_n8069_ & new_n8071_;
  assign new_n8073_ = ~new_n5105_ & new_n7990_;
  assign new_n8074_ = new_n8072_ & ~new_n8073_;
  assign new_n8075_ = new_n3815_ & new_n7985_;
  assign new_n8076_ = new_n4088_ & new_n7986_;
  assign new_n8077_ = ~new_n8075_ & ~new_n8076_;
  assign new_n8078_ = new_n3820_ & new_n7990_;
  assign new_n8079_ = new_n3870_ & new_n8036_;
  assign new_n8080_ = ~new_n8078_ & ~new_n8079_;
  assign new_n8081_ = ~new_n4069_ & new_n7986_;
  assign new_n8082_ = new_n8074_ & new_n8077_;
  assign new_n8083_ = new_n8080_ & new_n8082_;
  assign new_n8084_ = ~new_n8081_ & new_n8083_;
  assign new_n8085_ = new_n8064_ & new_n8084_;
  assign new_n8086_ = lo0062 & new_n5505_;
  assign new_n8087_ = lo0062 & new_n5135_;
  assign new_n8088_ = lo0062 & ~lo0993;
  assign new_n8089_ = new_n3927_ & new_n8088_;
  assign new_n8090_ = new_n3953_ & new_n7986_;
  assign new_n8091_ = ~new_n8089_ & ~new_n8090_;
  assign new_n8092_ = lo0024 & new_n4041_;
  assign new_n8093_ = ~new_n8086_ & ~new_n8087_;
  assign new_n8094_ = new_n8091_ & new_n8093_;
  assign new_n8095_ = ~new_n8092_ & new_n8094_;
  assign new_n8096_ = new_n8003_ & new_n8025_;
  assign new_n8097_ = new_n8085_ & new_n8096_;
  assign li0062 = ~new_n8095_ | ~new_n8097_;
  assign new_n8099_ = lo0063 & ~lo0314;
  assign new_n8100_ = ~lo0024 & lo0063;
  assign new_n8101_ = ~new_n5060_ & new_n8099_;
  assign new_n8102_ = new_n3940_ & new_n8100_;
  assign new_n8103_ = ~new_n8101_ & ~new_n8102_;
  assign new_n8104_ = lo0063 & ~lo0841;
  assign new_n8105_ = ~lo0024 & ~lo0063;
  assign new_n8106_ = lo0063 & new_n5194_;
  assign new_n8107_ = ~new_n8100_ & ~new_n8106_;
  assign new_n8108_ = new_n3936_ & ~new_n8107_;
  assign new_n8109_ = new_n3625_ & ~new_n8105_;
  assign new_n8110_ = ~new_n8108_ & ~new_n8109_;
  assign new_n8111_ = lo0063 & new_n3706_;
  assign new_n8112_ = lo0063 & new_n5818_;
  assign new_n8113_ = ~new_n5184_ & new_n8112_;
  assign new_n8114_ = new_n8110_ & ~new_n8111_;
  assign new_n8115_ = ~new_n8113_ & new_n8114_;
  assign new_n8116_ = ~new_n5201_ & new_n8104_;
  assign new_n8117_ = new_n8115_ & ~new_n8116_;
  assign new_n8118_ = new_n8103_ & new_n8117_;
  assign new_n8119_ = new_n4020_ & new_n8100_;
  assign new_n8120_ = ~new_n5096_ & new_n8104_;
  assign new_n8121_ = ~new_n8119_ & ~new_n8120_;
  assign new_n8122_ = lo0063 & new_n5071_;
  assign new_n8123_ = lo0063 & new_n4219_;
  assign new_n8124_ = lo0063 & li0583;
  assign new_n8125_ = ~new_n5074_ & new_n8123_;
  assign new_n8126_ = ~new_n5076_ & new_n8124_;
  assign new_n8127_ = ~new_n8125_ & ~new_n8126_;
  assign new_n8128_ = new_n4475_ & ~new_n8127_;
  assign new_n8129_ = lo0063 & new_n5083_;
  assign new_n8130_ = ~new_n8122_ & ~new_n8128_;
  assign new_n8131_ = ~new_n8129_ & new_n8130_;
  assign new_n8132_ = new_n5070_ & ~new_n8131_;
  assign new_n8133_ = ~new_n4096_ & new_n8100_;
  assign new_n8134_ = lo0063 & ~new_n8100_;
  assign new_n8135_ = ~new_n8133_ & ~new_n8134_;
  assign new_n8136_ = new_n5090_ & ~new_n8135_;
  assign new_n8137_ = new_n3746_ & new_n8099_;
  assign new_n8138_ = ~new_n8136_ & ~new_n8137_;
  assign new_n8139_ = new_n8121_ & ~new_n8132_;
  assign new_n8140_ = new_n8138_ & new_n8139_;
  assign new_n8141_ = lo0063 & ~new_n5216_;
  assign new_n8142_ = new_n4133_ & new_n8100_;
  assign new_n8143_ = ~new_n8141_ & ~new_n8142_;
  assign new_n8144_ = new_n3974_ & new_n8124_;
  assign new_n8145_ = ~new_n4135_ & new_n8144_;
  assign new_n8146_ = lo0063 & new_n5225_;
  assign new_n8147_ = new_n8143_ & ~new_n8145_;
  assign new_n8148_ = ~new_n8146_ & new_n8147_;
  assign new_n8149_ = new_n3948_ & new_n8100_;
  assign new_n8150_ = new_n8148_ & ~new_n8149_;
  assign new_n8151_ = lo0063 & new_n3678_;
  assign new_n8152_ = new_n3786_ & new_n8100_;
  assign new_n8153_ = new_n5139_ & new_n8151_;
  assign new_n8154_ = ~new_n8152_ & ~new_n8153_;
  assign new_n8155_ = new_n8150_ & new_n8154_;
  assign new_n8156_ = new_n4050_ & new_n8100_;
  assign new_n8157_ = lo0063 & new_n5562_;
  assign new_n8158_ = lo0063 & new_n5155_;
  assign new_n8159_ = new_n3777_ & new_n8158_;
  assign new_n8160_ = lo0063 & ~new_n4632_;
  assign new_n8161_ = new_n5565_ & new_n8160_;
  assign new_n8162_ = ~new_n8159_ & ~new_n8161_;
  assign new_n8163_ = ~new_n5460_ & new_n8099_;
  assign new_n8164_ = new_n8162_ & ~new_n8163_;
  assign new_n8165_ = new_n3763_ & new_n8104_;
  assign new_n8166_ = new_n3780_ & new_n8100_;
  assign new_n8167_ = ~new_n8165_ & ~new_n8166_;
  assign new_n8168_ = new_n3794_ & new_n8099_;
  assign new_n8169_ = new_n8167_ & ~new_n8168_;
  assign new_n8170_ = ~new_n8156_ & ~new_n8157_;
  assign new_n8171_ = new_n8164_ & new_n8170_;
  assign new_n8172_ = new_n8169_ & new_n8171_;
  assign new_n8173_ = new_n4041_ & new_n8100_;
  assign new_n8174_ = new_n8172_ & ~new_n8173_;
  assign new_n8175_ = new_n8155_ & new_n8174_;
  assign new_n8176_ = new_n3804_ & new_n8100_;
  assign new_n8177_ = new_n3834_ & new_n8124_;
  assign new_n8178_ = new_n3678_ & new_n8177_;
  assign new_n8179_ = lo0063 & new_n5112_;
  assign new_n8180_ = new_n3810_ & new_n8104_;
  assign new_n8181_ = ~new_n8176_ & ~new_n8178_;
  assign new_n8182_ = ~new_n8179_ & new_n8181_;
  assign new_n8183_ = ~new_n8180_ & new_n8182_;
  assign new_n8184_ = ~new_n5105_ & new_n8104_;
  assign new_n8185_ = new_n8183_ & ~new_n8184_;
  assign new_n8186_ = new_n3815_ & new_n8099_;
  assign new_n8187_ = new_n4088_ & new_n8100_;
  assign new_n8188_ = ~new_n8186_ & ~new_n8187_;
  assign new_n8189_ = ~lo1044 & new_n8099_;
  assign new_n8190_ = new_n3820_ & new_n8104_;
  assign new_n8191_ = new_n3870_ & new_n8189_;
  assign new_n8192_ = ~new_n8190_ & ~new_n8191_;
  assign new_n8193_ = ~new_n4069_ & new_n8100_;
  assign new_n8194_ = new_n8185_ & new_n8188_;
  assign new_n8195_ = new_n8192_ & new_n8194_;
  assign new_n8196_ = ~new_n8193_ & new_n8195_;
  assign new_n8197_ = new_n8175_ & new_n8196_;
  assign new_n8198_ = lo0063 & new_n5505_;
  assign new_n8199_ = lo0063 & new_n5135_;
  assign new_n8200_ = lo0063 & ~lo0993;
  assign new_n8201_ = new_n3927_ & new_n8200_;
  assign new_n8202_ = new_n3953_ & new_n8100_;
  assign new_n8203_ = ~new_n8201_ & ~new_n8202_;
  assign new_n8204_ = new_n4007_ & new_n8189_;
  assign new_n8205_ = new_n3969_ & new_n8104_;
  assign new_n8206_ = ~new_n8204_ & ~new_n8205_;
  assign new_n8207_ = ~new_n8198_ & ~new_n8199_;
  assign new_n8208_ = new_n8203_ & new_n8207_;
  assign new_n8209_ = new_n8206_ & new_n8208_;
  assign new_n8210_ = new_n8118_ & new_n8140_;
  assign new_n8211_ = new_n8197_ & new_n8210_;
  assign li0063 = ~new_n8209_ | ~new_n8211_;
  assign new_n8213_ = lo0064 & ~lo0314;
  assign new_n8214_ = ~lo0024 & lo0064;
  assign new_n8215_ = ~new_n5060_ & new_n8213_;
  assign new_n8216_ = new_n3940_ & new_n8214_;
  assign new_n8217_ = ~new_n8215_ & ~new_n8216_;
  assign new_n8218_ = lo0064 & ~lo0841;
  assign new_n8219_ = lo0064 & new_n5194_;
  assign new_n8220_ = ~new_n8214_ & ~new_n8219_;
  assign new_n8221_ = new_n3936_ & ~new_n8220_;
  assign new_n8222_ = new_n3625_ & new_n8214_;
  assign new_n8223_ = ~new_n8221_ & ~new_n8222_;
  assign new_n8224_ = lo0064 & new_n3706_;
  assign new_n8225_ = lo0064 & new_n5818_;
  assign new_n8226_ = ~new_n5184_ & new_n8225_;
  assign new_n8227_ = new_n8223_ & ~new_n8224_;
  assign new_n8228_ = ~new_n8226_ & new_n8227_;
  assign new_n8229_ = ~new_n5201_ & new_n8218_;
  assign new_n8230_ = new_n8228_ & ~new_n8229_;
  assign new_n8231_ = new_n8217_ & new_n8230_;
  assign new_n8232_ = new_n3804_ & new_n8214_;
  assign new_n8233_ = lo0064 & li0583;
  assign new_n8234_ = new_n3834_ & new_n8233_;
  assign new_n8235_ = new_n3678_ & new_n8234_;
  assign new_n8236_ = lo0064 & new_n5112_;
  assign new_n8237_ = new_n3810_ & new_n8218_;
  assign new_n8238_ = ~new_n8232_ & ~new_n8235_;
  assign new_n8239_ = ~new_n8236_ & new_n8238_;
  assign new_n8240_ = ~new_n8237_ & new_n8239_;
  assign new_n8241_ = ~new_n5105_ & new_n8218_;
  assign new_n8242_ = new_n8240_ & ~new_n8241_;
  assign new_n8243_ = new_n3815_ & new_n8213_;
  assign new_n8244_ = new_n4088_ & new_n8214_;
  assign new_n8245_ = ~new_n8243_ & ~new_n8244_;
  assign new_n8246_ = ~lo1044 & new_n8213_;
  assign new_n8247_ = new_n3820_ & new_n8218_;
  assign new_n8248_ = new_n3870_ & new_n8246_;
  assign new_n8249_ = ~new_n8247_ & ~new_n8248_;
  assign new_n8250_ = ~new_n4069_ & new_n8214_;
  assign new_n8251_ = new_n8242_ & new_n8245_;
  assign new_n8252_ = new_n8249_ & new_n8251_;
  assign new_n8253_ = ~new_n8250_ & new_n8252_;
  assign new_n8254_ = new_n3746_ & new_n8213_;
  assign new_n8255_ = new_n4020_ & new_n8214_;
  assign new_n8256_ = ~new_n8254_ & ~new_n8255_;
  assign new_n8257_ = ~new_n5096_ & new_n8218_;
  assign new_n8258_ = new_n8256_ & ~new_n8257_;
  assign new_n8259_ = lo0064 & new_n5071_;
  assign new_n8260_ = lo0064 & lo0786;
  assign new_n8261_ = ~new_n5076_ & new_n8233_;
  assign new_n8262_ = lo0064 & new_n5545_;
  assign new_n8263_ = ~new_n8261_ & ~new_n8262_;
  assign new_n8264_ = new_n4475_ & ~new_n8263_;
  assign new_n8265_ = new_n5082_ & new_n8260_;
  assign new_n8266_ = ~new_n8264_ & ~new_n8265_;
  assign new_n8267_ = ~new_n8259_ & new_n8266_;
  assign new_n8268_ = new_n4653_ & ~new_n8267_;
  assign new_n8269_ = ~new_n4096_ & new_n8214_;
  assign new_n8270_ = lo0064 & ~new_n8214_;
  assign new_n8271_ = ~new_n8269_ & ~new_n8270_;
  assign new_n8272_ = new_n4424_ & new_n8268_;
  assign new_n8273_ = new_n5090_ & ~new_n8271_;
  assign new_n8274_ = ~new_n8272_ & ~new_n8273_;
  assign new_n8275_ = new_n8258_ & new_n8274_;
  assign new_n8276_ = ~new_n3739_ & new_n8275_;
  assign new_n8277_ = new_n4050_ & new_n8214_;
  assign new_n8278_ = lo0064 & new_n5562_;
  assign new_n8279_ = lo0064 & new_n5155_;
  assign new_n8280_ = new_n3777_ & new_n8279_;
  assign new_n8281_ = lo0064 & ~new_n4632_;
  assign new_n8282_ = new_n5565_ & new_n8281_;
  assign new_n8283_ = ~new_n8280_ & ~new_n8282_;
  assign new_n8284_ = ~new_n5460_ & new_n8213_;
  assign new_n8285_ = new_n8283_ & ~new_n8284_;
  assign new_n8286_ = new_n3763_ & new_n8218_;
  assign new_n8287_ = new_n3780_ & new_n8214_;
  assign new_n8288_ = ~new_n8286_ & ~new_n8287_;
  assign new_n8289_ = new_n3794_ & new_n8213_;
  assign new_n8290_ = new_n8288_ & ~new_n8289_;
  assign new_n8291_ = ~new_n8277_ & ~new_n8278_;
  assign new_n8292_ = new_n8285_ & new_n8291_;
  assign new_n8293_ = new_n8290_ & new_n8292_;
  assign new_n8294_ = new_n4041_ & new_n8214_;
  assign new_n8295_ = new_n8293_ & ~new_n8294_;
  assign new_n8296_ = lo0064 & ~new_n5216_;
  assign new_n8297_ = new_n4133_ & new_n8214_;
  assign new_n8298_ = ~new_n8296_ & ~new_n8297_;
  assign new_n8299_ = new_n3974_ & new_n8233_;
  assign new_n8300_ = ~new_n4135_ & new_n8299_;
  assign new_n8301_ = lo0064 & new_n5225_;
  assign new_n8302_ = new_n8298_ & ~new_n8300_;
  assign new_n8303_ = ~new_n8301_ & new_n8302_;
  assign new_n8304_ = new_n3948_ & new_n8214_;
  assign new_n8305_ = new_n8303_ & ~new_n8304_;
  assign new_n8306_ = lo0064 & new_n3678_;
  assign new_n8307_ = new_n3786_ & new_n8214_;
  assign new_n8308_ = new_n5139_ & new_n8306_;
  assign new_n8309_ = ~new_n8307_ & ~new_n8308_;
  assign new_n8310_ = new_n8305_ & new_n8309_;
  assign new_n8311_ = new_n8295_ & new_n8310_;
  assign new_n8312_ = new_n8276_ & new_n8311_;
  assign new_n8313_ = lo0064 & new_n5505_;
  assign new_n8314_ = lo0064 & new_n5135_;
  assign new_n8315_ = lo0064 & ~lo0993;
  assign new_n8316_ = new_n3927_ & new_n8315_;
  assign new_n8317_ = new_n3953_ & new_n8214_;
  assign new_n8318_ = ~new_n8316_ & ~new_n8317_;
  assign new_n8319_ = new_n4007_ & new_n8246_;
  assign new_n8320_ = new_n3969_ & new_n8218_;
  assign new_n8321_ = ~new_n8319_ & ~new_n8320_;
  assign new_n8322_ = ~new_n8313_ & ~new_n8314_;
  assign new_n8323_ = new_n8318_ & new_n8322_;
  assign new_n8324_ = new_n8321_ & new_n8323_;
  assign new_n8325_ = new_n8231_ & new_n8253_;
  assign new_n8326_ = new_n8312_ & new_n8325_;
  assign li0064 = ~new_n8324_ | ~new_n8326_;
  assign new_n8328_ = ~lo0024 & lo0065;
  assign new_n8329_ = new_n4050_ & new_n8328_;
  assign new_n8330_ = lo0065 & new_n5562_;
  assign new_n8331_ = lo0065 & ~lo0314;
  assign new_n8332_ = lo0065 & new_n5155_;
  assign new_n8333_ = new_n3777_ & new_n8332_;
  assign new_n8334_ = lo0065 & ~new_n4632_;
  assign new_n8335_ = new_n5565_ & new_n8334_;
  assign new_n8336_ = ~new_n8333_ & ~new_n8335_;
  assign new_n8337_ = ~new_n5460_ & new_n8331_;
  assign new_n8338_ = new_n8336_ & ~new_n8337_;
  assign new_n8339_ = lo0065 & ~lo0841;
  assign new_n8340_ = new_n3763_ & new_n8339_;
  assign new_n8341_ = new_n3780_ & new_n8328_;
  assign new_n8342_ = ~new_n8340_ & ~new_n8341_;
  assign new_n8343_ = new_n3794_ & new_n8331_;
  assign new_n8344_ = new_n8342_ & ~new_n8343_;
  assign new_n8345_ = ~new_n8329_ & ~new_n8330_;
  assign new_n8346_ = new_n8338_ & new_n8345_;
  assign new_n8347_ = new_n8344_ & new_n8346_;
  assign new_n8348_ = new_n4041_ & new_n8328_;
  assign new_n8349_ = new_n8347_ & ~new_n8348_;
  assign new_n8350_ = lo0065 & ~new_n5216_;
  assign new_n8351_ = new_n4133_ & new_n8328_;
  assign new_n8352_ = ~new_n8350_ & ~new_n8351_;
  assign new_n8353_ = lo0065 & li0583;
  assign new_n8354_ = new_n3974_ & new_n8353_;
  assign new_n8355_ = ~new_n4135_ & new_n8354_;
  assign new_n8356_ = lo0065 & new_n5225_;
  assign new_n8357_ = new_n8352_ & ~new_n8355_;
  assign new_n8358_ = ~new_n8356_ & new_n8357_;
  assign new_n8359_ = new_n3948_ & new_n8328_;
  assign new_n8360_ = new_n8358_ & ~new_n8359_;
  assign new_n8361_ = lo0065 & new_n3678_;
  assign new_n8362_ = new_n3786_ & new_n8328_;
  assign new_n8363_ = new_n5139_ & new_n8361_;
  assign new_n8364_ = ~new_n8362_ & ~new_n8363_;
  assign new_n8365_ = new_n8360_ & new_n8364_;
  assign new_n8366_ = new_n8349_ & new_n8365_;
  assign new_n8367_ = new_n3804_ & new_n8328_;
  assign new_n8368_ = new_n3834_ & new_n8353_;
  assign new_n8369_ = new_n3678_ & new_n8368_;
  assign new_n8370_ = lo0065 & new_n5112_;
  assign new_n8371_ = new_n3810_ & new_n8339_;
  assign new_n8372_ = ~new_n8367_ & ~new_n8369_;
  assign new_n8373_ = ~new_n8370_ & new_n8372_;
  assign new_n8374_ = ~new_n8371_ & new_n8373_;
  assign new_n8375_ = ~new_n5105_ & new_n8339_;
  assign new_n8376_ = new_n8374_ & ~new_n8375_;
  assign new_n8377_ = new_n3815_ & new_n8331_;
  assign new_n8378_ = new_n4088_ & new_n8328_;
  assign new_n8379_ = ~new_n8377_ & ~new_n8378_;
  assign new_n8380_ = ~lo1044 & new_n8331_;
  assign new_n8381_ = new_n3820_ & new_n8339_;
  assign new_n8382_ = new_n3870_ & new_n8380_;
  assign new_n8383_ = ~new_n8381_ & ~new_n8382_;
  assign new_n8384_ = ~new_n4069_ & new_n8328_;
  assign new_n8385_ = new_n8376_ & new_n8379_;
  assign new_n8386_ = new_n8383_ & new_n8385_;
  assign new_n8387_ = ~new_n8384_ & new_n8386_;
  assign new_n8388_ = new_n8366_ & new_n8387_;
  assign new_n8389_ = lo0065 & new_n5505_;
  assign new_n8390_ = lo0065 & new_n5135_;
  assign new_n8391_ = lo0065 & ~lo0993;
  assign new_n8392_ = new_n3927_ & new_n8391_;
  assign new_n8393_ = new_n3953_ & new_n8328_;
  assign new_n8394_ = ~new_n8392_ & ~new_n8393_;
  assign new_n8395_ = new_n4007_ & new_n8380_;
  assign new_n8396_ = new_n3969_ & new_n8339_;
  assign new_n8397_ = ~new_n8395_ & ~new_n8396_;
  assign new_n8398_ = ~new_n8389_ & ~new_n8390_;
  assign new_n8399_ = new_n8394_ & new_n8398_;
  assign new_n8400_ = new_n8397_ & new_n8399_;
  assign new_n8401_ = new_n8388_ & new_n8400_;
  assign new_n8402_ = new_n4020_ & new_n8328_;
  assign new_n8403_ = ~new_n5096_ & new_n8339_;
  assign new_n8404_ = ~new_n8402_ & ~new_n8403_;
  assign new_n8405_ = lo0065 & new_n5071_;
  assign new_n8406_ = ~lo0065 & lo0786;
  assign new_n8407_ = ~new_n5076_ & new_n8353_;
  assign new_n8408_ = lo0065 & new_n5545_;
  assign new_n8409_ = ~new_n8407_ & ~new_n8408_;
  assign new_n8410_ = new_n4475_ & ~new_n8409_;
  assign new_n8411_ = new_n5082_ & ~new_n8406_;
  assign new_n8412_ = ~new_n8410_ & ~new_n8411_;
  assign new_n8413_ = ~new_n8405_ & new_n8412_;
  assign new_n8414_ = new_n5070_ & ~new_n8413_;
  assign new_n8415_ = ~new_n4096_ & new_n8328_;
  assign new_n8416_ = lo0065 & ~new_n8328_;
  assign new_n8417_ = ~new_n8415_ & ~new_n8416_;
  assign new_n8418_ = new_n5090_ & ~new_n8417_;
  assign new_n8419_ = new_n3746_ & new_n8331_;
  assign new_n8420_ = ~new_n8418_ & ~new_n8419_;
  assign new_n8421_ = new_n8404_ & ~new_n8414_;
  assign new_n8422_ = new_n8420_ & new_n8421_;
  assign new_n8423_ = ~new_n5060_ & new_n8331_;
  assign new_n8424_ = new_n3940_ & new_n8328_;
  assign new_n8425_ = ~new_n8423_ & ~new_n8424_;
  assign new_n8426_ = lo0065 & new_n5194_;
  assign new_n8427_ = ~new_n8328_ & ~new_n8426_;
  assign new_n8428_ = new_n3936_ & ~new_n8427_;
  assign new_n8429_ = new_n3625_ & new_n8328_;
  assign new_n8430_ = ~new_n8428_ & ~new_n8429_;
  assign new_n8431_ = lo0065 & new_n3706_;
  assign new_n8432_ = lo0065 & new_n5818_;
  assign new_n8433_ = ~new_n5184_ & new_n8432_;
  assign new_n8434_ = new_n8430_ & ~new_n8431_;
  assign new_n8435_ = ~new_n8433_ & new_n8434_;
  assign new_n8436_ = ~new_n5201_ & new_n8339_;
  assign new_n8437_ = new_n8435_ & ~new_n8436_;
  assign new_n8438_ = new_n8425_ & new_n8437_;
  assign new_n8439_ = new_n8422_ & new_n8438_;
  assign li0065 = ~new_n8401_ | ~new_n8439_;
  assign new_n8441_ = lo0066 & ~lo0314;
  assign new_n8442_ = ~lo0024 & lo0066;
  assign new_n8443_ = ~new_n5060_ & new_n8441_;
  assign new_n8444_ = new_n3940_ & new_n8442_;
  assign new_n8445_ = ~new_n8443_ & ~new_n8444_;
  assign new_n8446_ = lo0066 & ~lo0841;
  assign new_n8447_ = lo0066 & new_n5194_;
  assign new_n8448_ = ~new_n8442_ & ~new_n8447_;
  assign new_n8449_ = new_n3936_ & ~new_n8448_;
  assign new_n8450_ = new_n3625_ & new_n8442_;
  assign new_n8451_ = ~new_n8449_ & ~new_n8450_;
  assign new_n8452_ = lo0066 & new_n3706_;
  assign new_n8453_ = lo0066 & new_n5818_;
  assign new_n8454_ = ~new_n5184_ & new_n8453_;
  assign new_n8455_ = new_n8451_ & ~new_n8452_;
  assign new_n8456_ = ~new_n8454_ & new_n8455_;
  assign new_n8457_ = ~new_n5201_ & new_n8446_;
  assign new_n8458_ = new_n8456_ & ~new_n8457_;
  assign new_n8459_ = new_n8445_ & new_n8458_;
  assign new_n8460_ = new_n3804_ & new_n8442_;
  assign new_n8461_ = lo0066 & li0583;
  assign new_n8462_ = new_n3834_ & new_n8461_;
  assign new_n8463_ = new_n3678_ & new_n8462_;
  assign new_n8464_ = lo0066 & new_n5112_;
  assign new_n8465_ = new_n3810_ & new_n8446_;
  assign new_n8466_ = ~new_n8460_ & ~new_n8463_;
  assign new_n8467_ = ~new_n8464_ & new_n8466_;
  assign new_n8468_ = ~new_n8465_ & new_n8467_;
  assign new_n8469_ = ~new_n5105_ & new_n8446_;
  assign new_n8470_ = new_n8468_ & ~new_n8469_;
  assign new_n8471_ = new_n3815_ & new_n8441_;
  assign new_n8472_ = new_n4088_ & new_n8442_;
  assign new_n8473_ = ~new_n8471_ & ~new_n8472_;
  assign new_n8474_ = ~lo1044 & new_n8441_;
  assign new_n8475_ = new_n3820_ & new_n8446_;
  assign new_n8476_ = new_n3870_ & new_n8474_;
  assign new_n8477_ = ~new_n8475_ & ~new_n8476_;
  assign new_n8478_ = ~new_n4069_ & new_n8442_;
  assign new_n8479_ = new_n8470_ & new_n8473_;
  assign new_n8480_ = new_n8477_ & new_n8479_;
  assign new_n8481_ = ~new_n8478_ & new_n8480_;
  assign new_n8482_ = new_n4050_ & new_n8442_;
  assign new_n8483_ = lo0066 & new_n5562_;
  assign new_n8484_ = lo0066 & new_n5155_;
  assign new_n8485_ = new_n3777_ & new_n8484_;
  assign new_n8486_ = lo0066 & ~new_n4632_;
  assign new_n8487_ = new_n5565_ & new_n8486_;
  assign new_n8488_ = ~new_n8485_ & ~new_n8487_;
  assign new_n8489_ = ~new_n5460_ & new_n8441_;
  assign new_n8490_ = new_n8488_ & ~new_n8489_;
  assign new_n8491_ = new_n3763_ & new_n8446_;
  assign new_n8492_ = new_n3780_ & new_n8442_;
  assign new_n8493_ = ~new_n8491_ & ~new_n8492_;
  assign new_n8494_ = new_n3794_ & new_n8441_;
  assign new_n8495_ = new_n8493_ & ~new_n8494_;
  assign new_n8496_ = ~new_n8482_ & ~new_n8483_;
  assign new_n8497_ = new_n8490_ & new_n8496_;
  assign new_n8498_ = new_n8495_ & new_n8497_;
  assign new_n8499_ = new_n4041_ & new_n8442_;
  assign new_n8500_ = new_n8498_ & ~new_n8499_;
  assign new_n8501_ = lo0066 & ~new_n5216_;
  assign new_n8502_ = new_n4133_ & new_n8442_;
  assign new_n8503_ = ~new_n8501_ & ~new_n8502_;
  assign new_n8504_ = new_n3974_ & new_n8461_;
  assign new_n8505_ = ~new_n4135_ & new_n8504_;
  assign new_n8506_ = lo0066 & new_n5225_;
  assign new_n8507_ = new_n8503_ & ~new_n8505_;
  assign new_n8508_ = ~new_n8506_ & new_n8507_;
  assign new_n8509_ = new_n3948_ & new_n8442_;
  assign new_n8510_ = new_n8508_ & ~new_n8509_;
  assign new_n8511_ = lo0066 & new_n3678_;
  assign new_n8512_ = new_n3786_ & new_n8442_;
  assign new_n8513_ = new_n5139_ & new_n8511_;
  assign new_n8514_ = ~new_n8512_ & ~new_n8513_;
  assign new_n8515_ = new_n8510_ & new_n8514_;
  assign new_n8516_ = new_n8500_ & new_n8515_;
  assign new_n8517_ = new_n4020_ & new_n8442_;
  assign new_n8518_ = ~new_n5096_ & new_n8446_;
  assign new_n8519_ = ~new_n8517_ & ~new_n8518_;
  assign new_n8520_ = lo0066 & new_n5071_;
  assign new_n8521_ = lo0066 & lo0786;
  assign new_n8522_ = ~new_n5076_ & new_n8461_;
  assign new_n8523_ = lo0066 & new_n5545_;
  assign new_n8524_ = ~new_n8522_ & ~new_n8523_;
  assign new_n8525_ = new_n4475_ & ~new_n8524_;
  assign new_n8526_ = new_n5082_ & new_n8521_;
  assign new_n8527_ = ~new_n8525_ & ~new_n8526_;
  assign new_n8528_ = ~new_n8520_ & new_n8527_;
  assign new_n8529_ = new_n4653_ & ~new_n8528_;
  assign new_n8530_ = ~new_n4096_ & new_n8442_;
  assign new_n8531_ = lo0066 & ~new_n8442_;
  assign new_n8532_ = ~new_n8530_ & ~new_n8531_;
  assign new_n8533_ = new_n4424_ & new_n8529_;
  assign new_n8534_ = new_n5090_ & ~new_n8532_;
  assign new_n8535_ = ~new_n8533_ & ~new_n8534_;
  assign new_n8536_ = ~new_n6057_ & ~new_n6067_;
  assign new_n8537_ = lo0314 & ~new_n6074_;
  assign new_n8538_ = ~new_n8536_ & new_n8537_;
  assign new_n8539_ = ~new_n8441_ & ~new_n8538_;
  assign new_n8540_ = new_n3746_ & ~new_n8539_;
  assign new_n8541_ = new_n8519_ & new_n8535_;
  assign new_n8542_ = ~new_n8540_ & new_n8541_;
  assign new_n8543_ = new_n8516_ & new_n8542_;
  assign new_n8544_ = lo0066 & new_n5505_;
  assign new_n8545_ = lo0066 & new_n5135_;
  assign new_n8546_ = lo0066 & ~lo0993;
  assign new_n8547_ = new_n3927_ & new_n8546_;
  assign new_n8548_ = new_n3953_ & new_n8442_;
  assign new_n8549_ = ~new_n8547_ & ~new_n8548_;
  assign new_n8550_ = new_n4007_ & new_n8474_;
  assign new_n8551_ = new_n3969_ & new_n8446_;
  assign new_n8552_ = ~new_n8550_ & ~new_n8551_;
  assign new_n8553_ = ~new_n8544_ & ~new_n8545_;
  assign new_n8554_ = new_n8549_ & new_n8553_;
  assign new_n8555_ = new_n8552_ & new_n8554_;
  assign new_n8556_ = new_n8459_ & new_n8481_;
  assign new_n8557_ = new_n8543_ & new_n8556_;
  assign li0066 = ~new_n8555_ | ~new_n8557_;
  assign new_n8559_ = lo0067 & ~lo0314;
  assign new_n8560_ = ~lo0024 & lo0067;
  assign new_n8561_ = ~new_n5060_ & new_n8559_;
  assign new_n8562_ = new_n3940_ & new_n8560_;
  assign new_n8563_ = ~new_n8561_ & ~new_n8562_;
  assign new_n8564_ = lo0067 & ~lo0993;
  assign new_n8565_ = new_n3927_ & new_n8564_;
  assign new_n8566_ = new_n3953_ & new_n8560_;
  assign new_n8567_ = ~new_n8565_ & ~new_n8566_;
  assign new_n8568_ = new_n8563_ & new_n8567_;
  assign new_n8569_ = ~lo0067 & ~lo0314;
  assign new_n8570_ = new_n3903_ & ~new_n8569_;
  assign new_n8571_ = new_n3914_ & new_n8559_;
  assign new_n8572_ = ~new_n8570_ & ~new_n8571_;
  assign new_n8573_ = lo0067 & new_n6643_;
  assign new_n8574_ = lo0067 & ~new_n4632_;
  assign new_n8575_ = new_n5565_ & new_n8574_;
  assign new_n8576_ = new_n8572_ & ~new_n8573_;
  assign new_n8577_ = ~new_n8575_ & new_n8576_;
  assign new_n8578_ = new_n3794_ & new_n8559_;
  assign new_n8579_ = new_n8577_ & ~new_n8578_;
  assign new_n8580_ = lo0067 & new_n5562_;
  assign new_n8581_ = lo0067 & ~lo0841;
  assign new_n8582_ = new_n3780_ & new_n8560_;
  assign new_n8583_ = new_n3763_ & new_n8581_;
  assign new_n8584_ = ~new_n8582_ & ~new_n8583_;
  assign new_n8585_ = new_n4050_ & new_n8560_;
  assign new_n8586_ = new_n8579_ & ~new_n8580_;
  assign new_n8587_ = new_n8584_ & new_n8586_;
  assign new_n8588_ = ~new_n8585_ & new_n8587_;
  assign new_n8589_ = new_n4041_ & new_n8560_;
  assign new_n8590_ = new_n8588_ & ~new_n8589_;
  assign new_n8591_ = new_n3786_ & new_n8560_;
  assign new_n8592_ = lo0067 & new_n5140_;
  assign new_n8593_ = new_n8590_ & ~new_n8591_;
  assign new_n8594_ = ~new_n8592_ & new_n8593_;
  assign new_n8595_ = ~lo1044 & new_n8559_;
  assign new_n8596_ = new_n4007_ & new_n8595_;
  assign new_n8597_ = new_n3969_ & new_n8581_;
  assign new_n8598_ = ~new_n8596_ & ~new_n8597_;
  assign new_n8599_ = new_n3948_ & new_n8560_;
  assign new_n8600_ = lo0067 & li0583;
  assign new_n8601_ = new_n3974_ & new_n8600_;
  assign new_n8602_ = ~new_n4135_ & new_n8601_;
  assign new_n8603_ = lo0067 & new_n5225_;
  assign new_n8604_ = ~new_n8602_ & ~new_n8603_;
  assign new_n8605_ = lo0067 & ~new_n5216_;
  assign new_n8606_ = new_n4133_ & new_n8560_;
  assign new_n8607_ = ~new_n8605_ & ~new_n8606_;
  assign new_n8608_ = new_n8598_ & ~new_n8599_;
  assign new_n8609_ = new_n8604_ & new_n8608_;
  assign new_n8610_ = new_n8607_ & new_n8609_;
  assign new_n8611_ = new_n8594_ & new_n8610_;
  assign new_n8612_ = lo0067 & ~new_n5134_;
  assign new_n8613_ = ~new_n5201_ & new_n8581_;
  assign new_n8614_ = lo0067 & new_n5194_;
  assign new_n8615_ = ~new_n8560_ & ~new_n8614_;
  assign new_n8616_ = new_n3936_ & ~new_n8615_;
  assign new_n8617_ = new_n3625_ & new_n8560_;
  assign new_n8618_ = ~new_n8616_ & ~new_n8617_;
  assign new_n8619_ = lo0067 & new_n5608_;
  assign new_n8620_ = ~new_n5184_ & new_n8619_;
  assign new_n8621_ = lo0067 & new_n3706_;
  assign new_n8622_ = ~new_n8613_ & new_n8618_;
  assign new_n8623_ = ~new_n8620_ & new_n8622_;
  assign new_n8624_ = ~new_n8621_ & new_n8623_;
  assign new_n8625_ = new_n5133_ & new_n8612_;
  assign new_n8626_ = new_n8624_ & ~new_n8625_;
  assign new_n8627_ = lo0067 & new_n5505_;
  assign new_n8628_ = new_n8568_ & new_n8611_;
  assign new_n8629_ = new_n8626_ & new_n8628_;
  assign new_n8630_ = ~new_n8627_ & new_n8629_;
  assign new_n8631_ = new_n3804_ & new_n8560_;
  assign new_n8632_ = new_n3834_ & new_n8600_;
  assign new_n8633_ = new_n3678_ & new_n8632_;
  assign new_n8634_ = lo0067 & new_n5112_;
  assign new_n8635_ = new_n3810_ & new_n8581_;
  assign new_n8636_ = ~new_n8631_ & ~new_n8633_;
  assign new_n8637_ = ~new_n8634_ & new_n8636_;
  assign new_n8638_ = ~new_n8635_ & new_n8637_;
  assign new_n8639_ = ~new_n5105_ & new_n8581_;
  assign new_n8640_ = new_n8638_ & ~new_n8639_;
  assign new_n8641_ = new_n3815_ & new_n8559_;
  assign new_n8642_ = new_n4088_ & new_n8560_;
  assign new_n8643_ = ~new_n8641_ & ~new_n8642_;
  assign new_n8644_ = new_n3820_ & new_n8581_;
  assign new_n8645_ = new_n3870_ & new_n8595_;
  assign new_n8646_ = ~new_n8644_ & ~new_n8645_;
  assign new_n8647_ = ~new_n4069_ & new_n8560_;
  assign new_n8648_ = new_n8640_ & new_n8643_;
  assign new_n8649_ = new_n8646_ & new_n8648_;
  assign new_n8650_ = ~new_n8647_ & new_n8649_;
  assign new_n8651_ = new_n4020_ & new_n8560_;
  assign new_n8652_ = ~new_n5096_ & new_n8581_;
  assign new_n8653_ = ~new_n8651_ & ~new_n8652_;
  assign new_n8654_ = ~new_n4096_ & new_n8560_;
  assign new_n8655_ = lo0067 & ~new_n8560_;
  assign new_n8656_ = ~new_n8654_ & ~new_n8655_;
  assign new_n8657_ = new_n5090_ & ~new_n8656_;
  assign new_n8658_ = new_n3746_ & new_n8559_;
  assign new_n8659_ = ~new_n8657_ & ~new_n8658_;
  assign new_n8660_ = lo0067 & new_n5071_;
  assign new_n8661_ = lo0067 & new_n4219_;
  assign new_n8662_ = ~new_n5074_ & new_n8661_;
  assign new_n8663_ = ~new_n5076_ & new_n8600_;
  assign new_n8664_ = ~new_n8662_ & ~new_n8663_;
  assign new_n8665_ = new_n4475_ & ~new_n8664_;
  assign new_n8666_ = lo0067 & new_n5083_;
  assign new_n8667_ = ~new_n8660_ & ~new_n8665_;
  assign new_n8668_ = ~new_n8666_ & new_n8667_;
  assign new_n8669_ = new_n5070_ & ~new_n8668_;
  assign new_n8670_ = new_n8650_ & new_n8653_;
  assign new_n8671_ = new_n8659_ & new_n8670_;
  assign new_n8672_ = ~new_n8669_ & new_n8671_;
  assign li0067 = ~new_n8630_ | ~new_n8672_;
  assign new_n8674_ = ~lo0024 & lo0068;
  assign new_n8675_ = new_n4050_ & new_n8674_;
  assign new_n8676_ = lo0068 & new_n5562_;
  assign new_n8677_ = lo0068 & ~lo0314;
  assign new_n8678_ = lo0068 & new_n5155_;
  assign new_n8679_ = new_n3777_ & new_n8678_;
  assign new_n8680_ = lo0068 & ~new_n4632_;
  assign new_n8681_ = new_n5565_ & new_n8680_;
  assign new_n8682_ = ~new_n8679_ & ~new_n8681_;
  assign new_n8683_ = ~new_n5460_ & new_n8677_;
  assign new_n8684_ = new_n8682_ & ~new_n8683_;
  assign new_n8685_ = lo0068 & ~lo0841;
  assign new_n8686_ = new_n3763_ & new_n8685_;
  assign new_n8687_ = new_n3780_ & new_n8674_;
  assign new_n8688_ = ~new_n8686_ & ~new_n8687_;
  assign new_n8689_ = new_n3794_ & new_n8677_;
  assign new_n8690_ = new_n8688_ & ~new_n8689_;
  assign new_n8691_ = ~new_n8675_ & ~new_n8676_;
  assign new_n8692_ = new_n8684_ & new_n8691_;
  assign new_n8693_ = new_n8690_ & new_n8692_;
  assign new_n8694_ = new_n4041_ & new_n8674_;
  assign new_n8695_ = new_n8693_ & ~new_n8694_;
  assign new_n8696_ = lo0068 & ~new_n5216_;
  assign new_n8697_ = new_n4133_ & new_n8674_;
  assign new_n8698_ = ~new_n8696_ & ~new_n8697_;
  assign new_n8699_ = lo0068 & li0583;
  assign new_n8700_ = new_n3974_ & new_n8699_;
  assign new_n8701_ = ~new_n4135_ & new_n8700_;
  assign new_n8702_ = lo0068 & new_n5225_;
  assign new_n8703_ = new_n8698_ & ~new_n8701_;
  assign new_n8704_ = ~new_n8702_ & new_n8703_;
  assign new_n8705_ = new_n3948_ & new_n8674_;
  assign new_n8706_ = new_n8704_ & ~new_n8705_;
  assign new_n8707_ = lo0068 & new_n3678_;
  assign new_n8708_ = new_n3786_ & new_n8674_;
  assign new_n8709_ = new_n5139_ & new_n8707_;
  assign new_n8710_ = ~new_n8708_ & ~new_n8709_;
  assign new_n8711_ = new_n8706_ & new_n8710_;
  assign new_n8712_ = new_n8695_ & new_n8711_;
  assign new_n8713_ = new_n3804_ & new_n8674_;
  assign new_n8714_ = new_n3834_ & new_n8699_;
  assign new_n8715_ = new_n3678_ & new_n8714_;
  assign new_n8716_ = lo0068 & new_n5112_;
  assign new_n8717_ = new_n3810_ & new_n8685_;
  assign new_n8718_ = ~new_n8713_ & ~new_n8715_;
  assign new_n8719_ = ~new_n8716_ & new_n8718_;
  assign new_n8720_ = ~new_n8717_ & new_n8719_;
  assign new_n8721_ = ~new_n5105_ & new_n8685_;
  assign new_n8722_ = new_n8720_ & ~new_n8721_;
  assign new_n8723_ = new_n3815_ & new_n8677_;
  assign new_n8724_ = new_n4088_ & new_n8674_;
  assign new_n8725_ = ~new_n8723_ & ~new_n8724_;
  assign new_n8726_ = ~lo1044 & new_n8677_;
  assign new_n8727_ = new_n3820_ & new_n8685_;
  assign new_n8728_ = new_n3870_ & new_n8726_;
  assign new_n8729_ = ~new_n8727_ & ~new_n8728_;
  assign new_n8730_ = ~new_n4069_ & new_n8674_;
  assign new_n8731_ = new_n8722_ & new_n8725_;
  assign new_n8732_ = new_n8729_ & new_n8731_;
  assign new_n8733_ = ~new_n8730_ & new_n8732_;
  assign new_n8734_ = new_n8712_ & new_n8733_;
  assign new_n8735_ = lo0068 & new_n5505_;
  assign new_n8736_ = lo0068 & new_n5135_;
  assign new_n8737_ = lo0068 & ~lo0993;
  assign new_n8738_ = new_n3927_ & new_n8737_;
  assign new_n8739_ = new_n3953_ & new_n8674_;
  assign new_n8740_ = ~new_n8738_ & ~new_n8739_;
  assign new_n8741_ = new_n4007_ & new_n8726_;
  assign new_n8742_ = new_n3969_ & new_n8685_;
  assign new_n8743_ = ~new_n8741_ & ~new_n8742_;
  assign new_n8744_ = ~new_n8735_ & ~new_n8736_;
  assign new_n8745_ = new_n8740_ & new_n8744_;
  assign new_n8746_ = new_n8743_ & new_n8745_;
  assign new_n8747_ = new_n8734_ & new_n8746_;
  assign new_n8748_ = new_n4020_ & new_n8674_;
  assign new_n8749_ = ~new_n5096_ & new_n8685_;
  assign new_n8750_ = ~new_n8748_ & ~new_n8749_;
  assign new_n8751_ = lo0068 & new_n5071_;
  assign new_n8752_ = lo0068 & lo0786;
  assign new_n8753_ = lo0068 & new_n5545_;
  assign new_n8754_ = ~new_n5076_ & new_n8699_;
  assign new_n8755_ = new_n4228_ & new_n4528_;
  assign new_n8756_ = ~new_n8754_ & ~new_n8755_;
  assign new_n8757_ = ~new_n8753_ & new_n8756_;
  assign new_n8758_ = new_n4475_ & ~new_n8757_;
  assign new_n8759_ = new_n5082_ & new_n8752_;
  assign new_n8760_ = ~new_n8758_ & ~new_n8759_;
  assign new_n8761_ = ~new_n8751_ & new_n8760_;
  assign new_n8762_ = new_n5070_ & ~new_n8761_;
  assign new_n8763_ = ~new_n4096_ & new_n8674_;
  assign new_n8764_ = lo0068 & ~new_n8674_;
  assign new_n8765_ = ~new_n8763_ & ~new_n8764_;
  assign new_n8766_ = new_n5090_ & ~new_n8765_;
  assign new_n8767_ = new_n3746_ & new_n8677_;
  assign new_n8768_ = ~new_n8766_ & ~new_n8767_;
  assign new_n8769_ = new_n8750_ & ~new_n8762_;
  assign new_n8770_ = new_n8768_ & new_n8769_;
  assign new_n8771_ = ~new_n5060_ & new_n8677_;
  assign new_n8772_ = new_n3940_ & new_n8674_;
  assign new_n8773_ = ~new_n8771_ & ~new_n8772_;
  assign new_n8774_ = lo0068 & new_n5194_;
  assign new_n8775_ = ~new_n8674_ & ~new_n8774_;
  assign new_n8776_ = new_n3936_ & ~new_n8775_;
  assign new_n8777_ = new_n3625_ & new_n8674_;
  assign new_n8778_ = ~new_n8776_ & ~new_n8777_;
  assign new_n8779_ = lo0068 & new_n3706_;
  assign new_n8780_ = lo0068 & new_n5818_;
  assign new_n8781_ = ~new_n5184_ & new_n8780_;
  assign new_n8782_ = new_n8778_ & ~new_n8779_;
  assign new_n8783_ = ~new_n8781_ & new_n8782_;
  assign new_n8784_ = ~new_n5201_ & new_n8685_;
  assign new_n8785_ = new_n8783_ & ~new_n8784_;
  assign new_n8786_ = new_n8773_ & new_n8785_;
  assign new_n8787_ = new_n8770_ & new_n8786_;
  assign li0068 = ~new_n8747_ | ~new_n8787_;
  assign new_n8789_ = lo0069 & ~lo0841;
  assign new_n8790_ = ~new_n5201_ & new_n8789_;
  assign new_n8791_ = ~lo0024 & lo0069;
  assign new_n8792_ = lo0069 & new_n5194_;
  assign new_n8793_ = ~new_n8791_ & ~new_n8792_;
  assign new_n8794_ = new_n3936_ & ~new_n8793_;
  assign new_n8795_ = new_n3625_ & new_n8791_;
  assign new_n8796_ = ~new_n8794_ & ~new_n8795_;
  assign new_n8797_ = lo0069 & new_n5608_;
  assign new_n8798_ = ~new_n5184_ & new_n8797_;
  assign new_n8799_ = lo0069 & new_n3706_;
  assign new_n8800_ = ~new_n8790_ & new_n8796_;
  assign new_n8801_ = ~new_n8798_ & new_n8800_;
  assign new_n8802_ = ~new_n8799_ & new_n8801_;
  assign new_n8803_ = lo0069 & new_n5505_;
  assign new_n8804_ = lo0069 & ~lo0314;
  assign new_n8805_ = ~new_n5060_ & new_n8804_;
  assign new_n8806_ = new_n3940_ & new_n8791_;
  assign new_n8807_ = ~new_n8805_ & ~new_n8806_;
  assign new_n8808_ = lo0069 & ~lo0993;
  assign new_n8809_ = new_n3927_ & new_n8808_;
  assign new_n8810_ = new_n3953_ & new_n8791_;
  assign new_n8811_ = ~new_n8809_ & ~new_n8810_;
  assign new_n8812_ = new_n8807_ & new_n8811_;
  assign new_n8813_ = lo0069 & ~new_n5216_;
  assign new_n8814_ = new_n4133_ & new_n8791_;
  assign new_n8815_ = ~new_n8813_ & ~new_n8814_;
  assign new_n8816_ = ~lo1044 & new_n8804_;
  assign new_n8817_ = new_n4007_ & new_n8816_;
  assign new_n8818_ = new_n3969_ & new_n8789_;
  assign new_n8819_ = ~new_n8817_ & ~new_n8818_;
  assign new_n8820_ = new_n3948_ & new_n8791_;
  assign new_n8821_ = new_n8815_ & new_n8819_;
  assign new_n8822_ = ~new_n8820_ & new_n8821_;
  assign new_n8823_ = new_n8812_ & new_n8822_;
  assign new_n8824_ = lo0069 & li0583;
  assign new_n8825_ = new_n3974_ & new_n8824_;
  assign new_n8826_ = ~new_n4135_ & new_n8825_;
  assign new_n8827_ = lo0069 & new_n5225_;
  assign new_n8828_ = ~new_n8826_ & ~new_n8827_;
  assign new_n8829_ = ~new_n8803_ & new_n8823_;
  assign new_n8830_ = new_n8828_ & new_n8829_;
  assign new_n8831_ = new_n8802_ & new_n8830_;
  assign new_n8832_ = lo0069 & ~new_n5134_;
  assign new_n8833_ = lo0069 & new_n5562_;
  assign new_n8834_ = new_n4050_ & new_n8791_;
  assign new_n8835_ = ~new_n8833_ & ~new_n8834_;
  assign new_n8836_ = ~new_n4575_ & new_n8804_;
  assign new_n8837_ = new_n8835_ & ~new_n8836_;
  assign new_n8838_ = new_n3780_ & new_n8791_;
  assign new_n8839_ = new_n3763_ & new_n8789_;
  assign new_n8840_ = ~new_n8838_ & ~new_n8839_;
  assign new_n8841_ = lo0069 & new_n5155_;
  assign new_n8842_ = lo0069 & ~new_n4632_;
  assign new_n8843_ = new_n5565_ & new_n8842_;
  assign new_n8844_ = new_n3777_ & new_n8841_;
  assign new_n8845_ = ~new_n8843_ & ~new_n8844_;
  assign new_n8846_ = new_n3903_ & new_n8804_;
  assign new_n8847_ = ~new_n3907_ & ~new_n8846_;
  assign new_n8848_ = new_n8837_ & new_n8840_;
  assign new_n8849_ = new_n8845_ & new_n8848_;
  assign new_n8850_ = new_n8847_ & new_n8849_;
  assign new_n8851_ = new_n4041_ & new_n8791_;
  assign new_n8852_ = new_n8850_ & ~new_n8851_;
  assign new_n8853_ = new_n3786_ & new_n8791_;
  assign new_n8854_ = lo0069 & new_n5140_;
  assign new_n8855_ = new_n8852_ & ~new_n8853_;
  assign new_n8856_ = ~new_n8854_ & new_n8855_;
  assign new_n8857_ = new_n5133_ & new_n8832_;
  assign new_n8858_ = new_n8856_ & ~new_n8857_;
  assign new_n8859_ = new_n8831_ & new_n8858_;
  assign new_n8860_ = new_n3804_ & new_n8791_;
  assign new_n8861_ = new_n3834_ & new_n8824_;
  assign new_n8862_ = new_n3678_ & new_n8861_;
  assign new_n8863_ = lo0069 & new_n5112_;
  assign new_n8864_ = new_n3810_ & new_n8789_;
  assign new_n8865_ = ~new_n8860_ & ~new_n8862_;
  assign new_n8866_ = ~new_n8863_ & new_n8865_;
  assign new_n8867_ = ~new_n8864_ & new_n8866_;
  assign new_n8868_ = ~new_n5105_ & new_n8789_;
  assign new_n8869_ = new_n8867_ & ~new_n8868_;
  assign new_n8870_ = new_n3815_ & new_n8804_;
  assign new_n8871_ = new_n4088_ & new_n8791_;
  assign new_n8872_ = ~new_n8870_ & ~new_n8871_;
  assign new_n8873_ = new_n3820_ & new_n8789_;
  assign new_n8874_ = new_n3870_ & new_n8816_;
  assign new_n8875_ = ~new_n8873_ & ~new_n8874_;
  assign new_n8876_ = ~new_n4069_ & new_n8791_;
  assign new_n8877_ = new_n8869_ & new_n8872_;
  assign new_n8878_ = new_n8875_ & new_n8877_;
  assign new_n8879_ = ~new_n8876_ & new_n8878_;
  assign new_n8880_ = new_n4020_ & new_n8791_;
  assign new_n8881_ = ~new_n5096_ & new_n8789_;
  assign new_n8882_ = ~new_n8880_ & ~new_n8881_;
  assign new_n8883_ = ~new_n4096_ & new_n8791_;
  assign new_n8884_ = lo0069 & ~new_n8791_;
  assign new_n8885_ = ~new_n8883_ & ~new_n8884_;
  assign new_n8886_ = new_n5090_ & ~new_n8885_;
  assign new_n8887_ = new_n3746_ & new_n8804_;
  assign new_n8888_ = ~new_n8886_ & ~new_n8887_;
  assign new_n8889_ = lo0069 & new_n5071_;
  assign new_n8890_ = lo0069 & new_n4219_;
  assign new_n8891_ = ~new_n5074_ & new_n8890_;
  assign new_n8892_ = ~new_n5076_ & new_n8824_;
  assign new_n8893_ = ~new_n8891_ & ~new_n8892_;
  assign new_n8894_ = new_n4475_ & ~new_n8893_;
  assign new_n8895_ = lo0069 & new_n5083_;
  assign new_n8896_ = ~new_n8889_ & ~new_n8894_;
  assign new_n8897_ = ~new_n8895_ & new_n8896_;
  assign new_n8898_ = new_n5070_ & ~new_n8897_;
  assign new_n8899_ = new_n8879_ & new_n8882_;
  assign new_n8900_ = new_n8888_ & new_n8899_;
  assign new_n8901_ = ~new_n8898_ & new_n8900_;
  assign li0069 = ~new_n8859_ | ~new_n8901_;
  assign new_n8903_ = lo0070 & ~lo0841;
  assign new_n8904_ = ~lo0024 & lo0070;
  assign new_n8905_ = lo0070 & new_n5194_;
  assign new_n8906_ = ~new_n8904_ & ~new_n8905_;
  assign new_n8907_ = new_n3936_ & ~new_n8906_;
  assign new_n8908_ = new_n3625_ & new_n8904_;
  assign new_n8909_ = ~new_n8907_ & ~new_n8908_;
  assign new_n8910_ = lo0070 & new_n3706_;
  assign new_n8911_ = lo0070 & new_n5818_;
  assign new_n8912_ = ~new_n5184_ & new_n8911_;
  assign new_n8913_ = new_n8909_ & ~new_n8910_;
  assign new_n8914_ = ~new_n8912_ & new_n8913_;
  assign new_n8915_ = ~new_n5201_ & new_n8903_;
  assign new_n8916_ = new_n8914_ & ~new_n8915_;
  assign new_n8917_ = lo0070 & ~lo0314;
  assign new_n8918_ = ~new_n5060_ & new_n8917_;
  assign new_n8919_ = new_n3940_ & new_n8904_;
  assign new_n8920_ = ~new_n8918_ & ~new_n8919_;
  assign new_n8921_ = lo0070 & ~lo0993;
  assign new_n8922_ = new_n3927_ & new_n8921_;
  assign new_n8923_ = new_n3953_ & new_n8904_;
  assign new_n8924_ = ~new_n8922_ & ~new_n8923_;
  assign new_n8925_ = new_n8916_ & new_n8920_;
  assign new_n8926_ = new_n8924_ & new_n8925_;
  assign new_n8927_ = new_n3804_ & new_n8904_;
  assign new_n8928_ = lo0070 & li0583;
  assign new_n8929_ = new_n3834_ & new_n8928_;
  assign new_n8930_ = new_n3678_ & new_n8929_;
  assign new_n8931_ = lo0070 & new_n5112_;
  assign new_n8932_ = new_n3810_ & new_n8903_;
  assign new_n8933_ = ~new_n8927_ & ~new_n8930_;
  assign new_n8934_ = ~new_n8931_ & new_n8933_;
  assign new_n8935_ = ~new_n8932_ & new_n8934_;
  assign new_n8936_ = ~new_n5105_ & new_n8903_;
  assign new_n8937_ = new_n8935_ & ~new_n8936_;
  assign new_n8938_ = new_n3815_ & new_n8917_;
  assign new_n8939_ = new_n4088_ & new_n8904_;
  assign new_n8940_ = ~new_n8938_ & ~new_n8939_;
  assign new_n8941_ = ~lo1044 & new_n8917_;
  assign new_n8942_ = new_n3820_ & new_n8903_;
  assign new_n8943_ = new_n3870_ & new_n8941_;
  assign new_n8944_ = ~new_n8942_ & ~new_n8943_;
  assign new_n8945_ = ~new_n4069_ & new_n8904_;
  assign new_n8946_ = new_n8937_ & new_n8940_;
  assign new_n8947_ = new_n8944_ & new_n8946_;
  assign new_n8948_ = ~new_n8945_ & new_n8947_;
  assign new_n8949_ = new_n4020_ & new_n8904_;
  assign new_n8950_ = ~new_n5096_ & new_n8903_;
  assign new_n8951_ = ~new_n8949_ & ~new_n8950_;
  assign new_n8952_ = ~new_n4096_ & new_n8904_;
  assign new_n8953_ = lo0070 & ~new_n8904_;
  assign new_n8954_ = ~new_n8952_ & ~new_n8953_;
  assign new_n8955_ = new_n5090_ & ~new_n8954_;
  assign new_n8956_ = new_n3746_ & new_n8917_;
  assign new_n8957_ = ~new_n8955_ & ~new_n8956_;
  assign new_n8958_ = lo0070 & new_n5071_;
  assign new_n8959_ = lo0070 & new_n5083_;
  assign new_n8960_ = lo0589 & ~new_n4053_;
  assign new_n8961_ = lo0593 & new_n8960_;
  assign new_n8962_ = new_n8960_ & ~new_n8961_;
  assign new_n8963_ = new_n5074_ & ~new_n8962_;
  assign new_n8964_ = ~lo0070 & ~new_n5074_;
  assign new_n8965_ = ~new_n8963_ & ~new_n8964_;
  assign new_n8966_ = new_n4219_ & new_n8965_;
  assign new_n8967_ = ~new_n5076_ & new_n8928_;
  assign new_n8968_ = ~new_n8966_ & ~new_n8967_;
  assign new_n8969_ = new_n4475_ & ~new_n8968_;
  assign new_n8970_ = ~new_n8958_ & ~new_n8959_;
  assign new_n8971_ = ~new_n8969_ & new_n8970_;
  assign new_n8972_ = new_n3612_ & ~new_n8971_;
  assign new_n8973_ = new_n4424_ & new_n8972_;
  assign new_n8974_ = ~new_n4482_ & new_n8951_;
  assign new_n8975_ = new_n8957_ & new_n8974_;
  assign new_n8976_ = ~new_n8973_ & new_n8975_;
  assign new_n8977_ = new_n8948_ & new_n8976_;
  assign new_n8978_ = lo0070 & new_n5505_;
  assign new_n8979_ = lo0070 & new_n5135_;
  assign new_n8980_ = new_n4007_ & new_n8941_;
  assign new_n8981_ = new_n3969_ & new_n8903_;
  assign new_n8982_ = ~new_n8980_ & ~new_n8981_;
  assign new_n8983_ = ~new_n8978_ & ~new_n8979_;
  assign new_n8984_ = new_n8982_ & new_n8983_;
  assign new_n8985_ = new_n4050_ & new_n8904_;
  assign new_n8986_ = lo0070 & new_n5562_;
  assign new_n8987_ = lo0070 & new_n5155_;
  assign new_n8988_ = new_n3777_ & new_n8987_;
  assign new_n8989_ = lo0070 & ~new_n4632_;
  assign new_n8990_ = new_n5565_ & new_n8989_;
  assign new_n8991_ = ~new_n8988_ & ~new_n8990_;
  assign new_n8992_ = ~new_n5460_ & new_n8917_;
  assign new_n8993_ = new_n8991_ & ~new_n8992_;
  assign new_n8994_ = new_n3763_ & new_n8903_;
  assign new_n8995_ = new_n3780_ & new_n8904_;
  assign new_n8996_ = ~new_n8994_ & ~new_n8995_;
  assign new_n8997_ = new_n3794_ & new_n8917_;
  assign new_n8998_ = new_n8996_ & ~new_n8997_;
  assign new_n8999_ = ~new_n8985_ & ~new_n8986_;
  assign new_n9000_ = new_n8993_ & new_n8999_;
  assign new_n9001_ = new_n8998_ & new_n9000_;
  assign new_n9002_ = new_n4041_ & new_n8904_;
  assign new_n9003_ = new_n9001_ & ~new_n9002_;
  assign new_n9004_ = lo0070 & ~new_n5216_;
  assign new_n9005_ = new_n4133_ & new_n8904_;
  assign new_n9006_ = ~new_n9004_ & ~new_n9005_;
  assign new_n9007_ = new_n3974_ & new_n8928_;
  assign new_n9008_ = ~new_n4135_ & new_n9007_;
  assign new_n9009_ = lo0070 & new_n5225_;
  assign new_n9010_ = new_n9006_ & ~new_n9008_;
  assign new_n9011_ = ~new_n9009_ & new_n9010_;
  assign new_n9012_ = new_n3948_ & new_n8904_;
  assign new_n9013_ = new_n9011_ & ~new_n9012_;
  assign new_n9014_ = lo0070 & new_n3678_;
  assign new_n9015_ = new_n3786_ & new_n8904_;
  assign new_n9016_ = new_n5139_ & new_n9014_;
  assign new_n9017_ = ~new_n9015_ & ~new_n9016_;
  assign new_n9018_ = new_n9003_ & new_n9013_;
  assign new_n9019_ = new_n9017_ & new_n9018_;
  assign new_n9020_ = new_n8984_ & new_n9019_;
  assign new_n9021_ = new_n8926_ & new_n8977_;
  assign li0070 = ~new_n9020_ | ~new_n9021_;
  assign new_n9023_ = lo0071 & new_n5505_;
  assign new_n9024_ = ~lo0024 & lo0071;
  assign new_n9025_ = lo0071 & ~lo0314;
  assign new_n9026_ = ~lo0071 & ~lo0314;
  assign new_n9027_ = new_n3914_ & ~new_n9026_;
  assign new_n9028_ = new_n3903_ & new_n9025_;
  assign new_n9029_ = ~new_n9027_ & ~new_n9028_;
  assign new_n9030_ = lo0071 & new_n6643_;
  assign new_n9031_ = lo0071 & ~new_n4632_;
  assign new_n9032_ = new_n5565_ & new_n9031_;
  assign new_n9033_ = new_n9029_ & ~new_n9030_;
  assign new_n9034_ = ~new_n9032_ & new_n9033_;
  assign new_n9035_ = new_n3794_ & new_n9025_;
  assign new_n9036_ = new_n9034_ & ~new_n9035_;
  assign new_n9037_ = lo0071 & new_n5562_;
  assign new_n9038_ = lo0071 & ~lo0841;
  assign new_n9039_ = new_n3780_ & new_n9024_;
  assign new_n9040_ = new_n3763_ & new_n9038_;
  assign new_n9041_ = ~new_n9039_ & ~new_n9040_;
  assign new_n9042_ = new_n4050_ & new_n9024_;
  assign new_n9043_ = new_n9036_ & ~new_n9037_;
  assign new_n9044_ = new_n9041_ & new_n9043_;
  assign new_n9045_ = ~new_n9042_ & new_n9044_;
  assign new_n9046_ = new_n4041_ & new_n9024_;
  assign new_n9047_ = new_n9045_ & ~new_n9046_;
  assign new_n9048_ = new_n3786_ & new_n9024_;
  assign new_n9049_ = lo0071 & new_n5140_;
  assign new_n9050_ = new_n9047_ & ~new_n9048_;
  assign new_n9051_ = ~new_n9049_ & new_n9050_;
  assign new_n9052_ = ~lo1044 & new_n9025_;
  assign new_n9053_ = new_n4007_ & new_n9052_;
  assign new_n9054_ = new_n3969_ & new_n9038_;
  assign new_n9055_ = ~new_n9053_ & ~new_n9054_;
  assign new_n9056_ = new_n3948_ & new_n9024_;
  assign new_n9057_ = lo0071 & li0583;
  assign new_n9058_ = new_n3974_ & new_n9057_;
  assign new_n9059_ = ~new_n4135_ & new_n9058_;
  assign new_n9060_ = lo0071 & new_n5225_;
  assign new_n9061_ = ~new_n9059_ & ~new_n9060_;
  assign new_n9062_ = lo0071 & ~new_n5216_;
  assign new_n9063_ = new_n4133_ & new_n9024_;
  assign new_n9064_ = ~new_n9062_ & ~new_n9063_;
  assign new_n9065_ = new_n9055_ & ~new_n9056_;
  assign new_n9066_ = new_n9061_ & new_n9065_;
  assign new_n9067_ = new_n9064_ & new_n9066_;
  assign new_n9068_ = new_n9051_ & new_n9067_;
  assign new_n9069_ = lo0071 & ~new_n5134_;
  assign new_n9070_ = ~new_n5201_ & new_n9038_;
  assign new_n9071_ = lo0071 & new_n5194_;
  assign new_n9072_ = ~new_n9024_ & ~new_n9071_;
  assign new_n9073_ = new_n3936_ & ~new_n9072_;
  assign new_n9074_ = new_n3625_ & new_n9024_;
  assign new_n9075_ = ~new_n9073_ & ~new_n9074_;
  assign new_n9076_ = lo0071 & new_n5608_;
  assign new_n9077_ = ~new_n5184_ & new_n9076_;
  assign new_n9078_ = lo0071 & new_n3706_;
  assign new_n9079_ = ~new_n9070_ & new_n9075_;
  assign new_n9080_ = ~new_n9077_ & new_n9079_;
  assign new_n9081_ = ~new_n9078_ & new_n9080_;
  assign new_n9082_ = new_n5133_ & new_n9069_;
  assign new_n9083_ = new_n9081_ & ~new_n9082_;
  assign new_n9084_ = ~new_n5060_ & new_n9025_;
  assign new_n9085_ = new_n3940_ & new_n9024_;
  assign new_n9086_ = ~new_n9084_ & ~new_n9085_;
  assign new_n9087_ = lo0071 & ~lo0993;
  assign new_n9088_ = new_n3927_ & new_n9087_;
  assign new_n9089_ = new_n3953_ & new_n9024_;
  assign new_n9090_ = ~new_n9088_ & ~new_n9089_;
  assign new_n9091_ = new_n9086_ & new_n9090_;
  assign new_n9092_ = ~new_n9023_ & new_n9068_;
  assign new_n9093_ = new_n9083_ & new_n9092_;
  assign new_n9094_ = new_n9091_ & new_n9093_;
  assign new_n9095_ = new_n3804_ & new_n9024_;
  assign new_n9096_ = new_n3834_ & new_n9057_;
  assign new_n9097_ = new_n3678_ & new_n9096_;
  assign new_n9098_ = lo0071 & new_n5112_;
  assign new_n9099_ = new_n3810_ & new_n9038_;
  assign new_n9100_ = ~new_n9095_ & ~new_n9097_;
  assign new_n9101_ = ~new_n9098_ & new_n9100_;
  assign new_n9102_ = ~new_n9099_ & new_n9101_;
  assign new_n9103_ = ~new_n5105_ & new_n9038_;
  assign new_n9104_ = new_n9102_ & ~new_n9103_;
  assign new_n9105_ = new_n3815_ & new_n9025_;
  assign new_n9106_ = new_n4088_ & new_n9024_;
  assign new_n9107_ = ~new_n9105_ & ~new_n9106_;
  assign new_n9108_ = new_n3820_ & new_n9038_;
  assign new_n9109_ = new_n3870_ & new_n9052_;
  assign new_n9110_ = ~new_n9108_ & ~new_n9109_;
  assign new_n9111_ = ~new_n4069_ & new_n9024_;
  assign new_n9112_ = new_n9104_ & new_n9107_;
  assign new_n9113_ = new_n9110_ & new_n9112_;
  assign new_n9114_ = ~new_n9111_ & new_n9113_;
  assign new_n9115_ = new_n4020_ & new_n9024_;
  assign new_n9116_ = ~new_n5096_ & new_n9038_;
  assign new_n9117_ = ~new_n9115_ & ~new_n9116_;
  assign new_n9118_ = new_n8536_ & new_n8537_;
  assign new_n9119_ = ~new_n9025_ & ~new_n9118_;
  assign new_n9120_ = new_n3746_ & ~new_n9119_;
  assign new_n9121_ = lo0071 & new_n5071_;
  assign new_n9122_ = lo0071 & lo0786;
  assign new_n9123_ = ~new_n5076_ & new_n9057_;
  assign new_n9124_ = lo0071 & new_n5545_;
  assign new_n9125_ = ~new_n9123_ & ~new_n9124_;
  assign new_n9126_ = new_n4475_ & ~new_n9125_;
  assign new_n9127_ = new_n5082_ & new_n9122_;
  assign new_n9128_ = ~new_n9126_ & ~new_n9127_;
  assign new_n9129_ = ~new_n9121_ & new_n9128_;
  assign new_n9130_ = new_n4653_ & ~new_n9129_;
  assign new_n9131_ = ~new_n4096_ & new_n9024_;
  assign new_n9132_ = lo0071 & ~new_n9024_;
  assign new_n9133_ = ~new_n9131_ & ~new_n9132_;
  assign new_n9134_ = new_n4424_ & new_n9130_;
  assign new_n9135_ = new_n5090_ & ~new_n9133_;
  assign new_n9136_ = ~new_n9134_ & ~new_n9135_;
  assign new_n9137_ = new_n9114_ & new_n9117_;
  assign new_n9138_ = ~new_n9120_ & new_n9137_;
  assign new_n9139_ = new_n9136_ & new_n9138_;
  assign li0071 = ~new_n9094_ | ~new_n9139_;
  assign new_n9141_ = lo0072 & ~lo0314;
  assign new_n9142_ = ~lo0024 & lo0072;
  assign new_n9143_ = ~new_n5060_ & new_n9141_;
  assign new_n9144_ = new_n3940_ & new_n9142_;
  assign new_n9145_ = ~new_n9143_ & ~new_n9144_;
  assign new_n9146_ = lo0072 & ~lo0993;
  assign new_n9147_ = new_n3927_ & new_n9146_;
  assign new_n9148_ = new_n3953_ & new_n9142_;
  assign new_n9149_ = ~new_n9147_ & ~new_n9148_;
  assign new_n9150_ = new_n9145_ & new_n9149_;
  assign new_n9151_ = new_n4050_ & new_n9142_;
  assign new_n9152_ = lo0072 & new_n5562_;
  assign new_n9153_ = lo0072 & new_n5155_;
  assign new_n9154_ = new_n3777_ & new_n9153_;
  assign new_n9155_ = lo0072 & ~new_n4632_;
  assign new_n9156_ = new_n5565_ & new_n9155_;
  assign new_n9157_ = ~new_n9154_ & ~new_n9156_;
  assign new_n9158_ = ~new_n5460_ & new_n9141_;
  assign new_n9159_ = new_n9157_ & ~new_n9158_;
  assign new_n9160_ = lo0072 & ~lo0841;
  assign new_n9161_ = new_n3763_ & new_n9160_;
  assign new_n9162_ = new_n3780_ & new_n9142_;
  assign new_n9163_ = ~new_n9161_ & ~new_n9162_;
  assign new_n9164_ = new_n3794_ & new_n9141_;
  assign new_n9165_ = new_n9163_ & ~new_n9164_;
  assign new_n9166_ = ~new_n9151_ & ~new_n9152_;
  assign new_n9167_ = new_n9159_ & new_n9166_;
  assign new_n9168_ = new_n9165_ & new_n9167_;
  assign new_n9169_ = new_n4041_ & new_n9142_;
  assign new_n9170_ = new_n9168_ & ~new_n9169_;
  assign new_n9171_ = lo0072 & new_n3678_;
  assign new_n9172_ = new_n3786_ & new_n9142_;
  assign new_n9173_ = new_n5139_ & new_n9171_;
  assign new_n9174_ = ~new_n9172_ & ~new_n9173_;
  assign new_n9175_ = ~lo1044 & new_n9141_;
  assign new_n9176_ = new_n4007_ & new_n9175_;
  assign new_n9177_ = new_n3969_ & new_n9160_;
  assign new_n9178_ = ~new_n9176_ & ~new_n9177_;
  assign new_n9179_ = lo0072 & ~new_n5216_;
  assign new_n9180_ = new_n4133_ & new_n9142_;
  assign new_n9181_ = ~new_n9179_ & ~new_n9180_;
  assign new_n9182_ = lo0072 & li0583;
  assign new_n9183_ = new_n3974_ & new_n9182_;
  assign new_n9184_ = ~new_n4135_ & new_n9183_;
  assign new_n9185_ = lo0072 & new_n5225_;
  assign new_n9186_ = new_n9181_ & ~new_n9184_;
  assign new_n9187_ = ~new_n9185_ & new_n9186_;
  assign new_n9188_ = new_n3948_ & new_n9142_;
  assign new_n9189_ = new_n9187_ & ~new_n9188_;
  assign new_n9190_ = new_n9170_ & new_n9174_;
  assign new_n9191_ = new_n9178_ & new_n9190_;
  assign new_n9192_ = new_n9189_ & new_n9191_;
  assign new_n9193_ = lo0072 & ~new_n5134_;
  assign new_n9194_ = ~new_n5201_ & new_n9160_;
  assign new_n9195_ = lo0072 & new_n5194_;
  assign new_n9196_ = ~new_n9142_ & ~new_n9195_;
  assign new_n9197_ = new_n3936_ & ~new_n9196_;
  assign new_n9198_ = new_n3625_ & new_n9142_;
  assign new_n9199_ = ~new_n9197_ & ~new_n9198_;
  assign new_n9200_ = lo0072 & new_n5708_;
  assign new_n9201_ = lo0072 & new_n3706_;
  assign new_n9202_ = ~new_n9194_ & new_n9199_;
  assign new_n9203_ = ~new_n9200_ & new_n9202_;
  assign new_n9204_ = ~new_n9201_ & new_n9203_;
  assign new_n9205_ = new_n5133_ & new_n9193_;
  assign new_n9206_ = new_n9204_ & ~new_n9205_;
  assign new_n9207_ = lo0072 & new_n5505_;
  assign new_n9208_ = new_n9150_ & new_n9192_;
  assign new_n9209_ = new_n9206_ & new_n9208_;
  assign new_n9210_ = ~new_n9207_ & new_n9209_;
  assign new_n9211_ = new_n3804_ & new_n9142_;
  assign new_n9212_ = new_n3834_ & new_n9171_;
  assign new_n9213_ = ~new_n9211_ & ~new_n9212_;
  assign new_n9214_ = ~li0583 & new_n3834_;
  assign new_n9215_ = new_n3678_ & new_n9214_;
  assign new_n9216_ = lo0072 & new_n5112_;
  assign new_n9217_ = new_n3810_ & new_n9160_;
  assign new_n9218_ = new_n9213_ & ~new_n9215_;
  assign new_n9219_ = ~new_n9216_ & new_n9218_;
  assign new_n9220_ = ~new_n9217_ & new_n9219_;
  assign new_n9221_ = ~new_n5105_ & new_n9160_;
  assign new_n9222_ = new_n9220_ & ~new_n9221_;
  assign new_n9223_ = new_n3815_ & new_n9141_;
  assign new_n9224_ = new_n4088_ & new_n9142_;
  assign new_n9225_ = ~new_n9223_ & ~new_n9224_;
  assign new_n9226_ = new_n3820_ & new_n9160_;
  assign new_n9227_ = new_n3870_ & new_n9175_;
  assign new_n9228_ = ~new_n9226_ & ~new_n9227_;
  assign new_n9229_ = ~new_n4069_ & new_n9142_;
  assign new_n9230_ = new_n9222_ & new_n9225_;
  assign new_n9231_ = new_n9228_ & new_n9230_;
  assign new_n9232_ = ~new_n9229_ & new_n9231_;
  assign new_n9233_ = new_n4020_ & new_n9142_;
  assign new_n9234_ = ~new_n5096_ & new_n9160_;
  assign new_n9235_ = ~new_n9233_ & ~new_n9234_;
  assign new_n9236_ = ~new_n4096_ & new_n9142_;
  assign new_n9237_ = lo0072 & ~new_n9142_;
  assign new_n9238_ = ~new_n9236_ & ~new_n9237_;
  assign new_n9239_ = new_n5090_ & ~new_n9238_;
  assign new_n9240_ = new_n3746_ & new_n9141_;
  assign new_n9241_ = ~new_n9239_ & ~new_n9240_;
  assign new_n9242_ = lo0072 & new_n5071_;
  assign new_n9243_ = lo0072 & lo0786;
  assign new_n9244_ = lo0072 & new_n5545_;
  assign new_n9245_ = ~new_n5076_ & new_n9182_;
  assign new_n9246_ = ~new_n4529_ & ~new_n9245_;
  assign new_n9247_ = ~new_n9244_ & new_n9246_;
  assign new_n9248_ = new_n4475_ & ~new_n9247_;
  assign new_n9249_ = new_n5082_ & new_n9243_;
  assign new_n9250_ = ~new_n9248_ & ~new_n9249_;
  assign new_n9251_ = ~new_n9242_ & new_n9250_;
  assign new_n9252_ = new_n5070_ & ~new_n9251_;
  assign new_n9253_ = new_n9232_ & new_n9235_;
  assign new_n9254_ = new_n9241_ & new_n9253_;
  assign new_n9255_ = ~new_n9252_ & new_n9254_;
  assign li0072 = ~new_n9210_ | ~new_n9255_;
  assign new_n9257_ = lo0073 & ~lo0314;
  assign new_n9258_ = ~lo0024 & lo0073;
  assign new_n9259_ = ~new_n5060_ & new_n9257_;
  assign new_n9260_ = new_n3940_ & new_n9258_;
  assign new_n9261_ = ~new_n9259_ & ~new_n9260_;
  assign new_n9262_ = lo0073 & ~lo0993;
  assign new_n9263_ = new_n3927_ & new_n9262_;
  assign new_n9264_ = new_n3953_ & new_n9258_;
  assign new_n9265_ = ~new_n9263_ & ~new_n9264_;
  assign new_n9266_ = new_n9261_ & new_n9265_;
  assign new_n9267_ = new_n4050_ & new_n9258_;
  assign new_n9268_ = lo0073 & new_n5562_;
  assign new_n9269_ = lo0073 & new_n5155_;
  assign new_n9270_ = new_n3777_ & new_n9269_;
  assign new_n9271_ = lo0073 & ~new_n4632_;
  assign new_n9272_ = new_n5565_ & new_n9271_;
  assign new_n9273_ = ~new_n9270_ & ~new_n9272_;
  assign new_n9274_ = ~new_n5460_ & new_n9257_;
  assign new_n9275_ = new_n9273_ & ~new_n9274_;
  assign new_n9276_ = lo0073 & ~lo0841;
  assign new_n9277_ = new_n3763_ & new_n9276_;
  assign new_n9278_ = new_n3780_ & new_n9258_;
  assign new_n9279_ = ~new_n9277_ & ~new_n9278_;
  assign new_n9280_ = new_n3794_ & new_n9257_;
  assign new_n9281_ = new_n9279_ & ~new_n9280_;
  assign new_n9282_ = ~new_n9267_ & ~new_n9268_;
  assign new_n9283_ = new_n9275_ & new_n9282_;
  assign new_n9284_ = new_n9281_ & new_n9283_;
  assign new_n9285_ = new_n4041_ & new_n9258_;
  assign new_n9286_ = new_n9284_ & ~new_n9285_;
  assign new_n9287_ = new_n3786_ & new_n9258_;
  assign new_n9288_ = lo0073 & new_n5140_;
  assign new_n9289_ = new_n9286_ & ~new_n9287_;
  assign new_n9290_ = ~new_n9288_ & new_n9289_;
  assign new_n9291_ = ~lo1044 & new_n9257_;
  assign new_n9292_ = new_n4007_ & new_n9291_;
  assign new_n9293_ = new_n3969_ & new_n9276_;
  assign new_n9294_ = ~new_n9292_ & ~new_n9293_;
  assign new_n9295_ = new_n3948_ & new_n9258_;
  assign new_n9296_ = lo0073 & li0583;
  assign new_n9297_ = new_n3974_ & new_n9296_;
  assign new_n9298_ = ~new_n4135_ & new_n9297_;
  assign new_n9299_ = lo0073 & new_n5225_;
  assign new_n9300_ = ~new_n9298_ & ~new_n9299_;
  assign new_n9301_ = lo0073 & ~new_n5216_;
  assign new_n9302_ = new_n4133_ & new_n9258_;
  assign new_n9303_ = ~new_n9301_ & ~new_n9302_;
  assign new_n9304_ = new_n9294_ & ~new_n9295_;
  assign new_n9305_ = new_n9300_ & new_n9304_;
  assign new_n9306_ = new_n9303_ & new_n9305_;
  assign new_n9307_ = new_n9290_ & new_n9306_;
  assign new_n9308_ = lo0073 & ~new_n5134_;
  assign new_n9309_ = ~new_n5201_ & new_n9276_;
  assign new_n9310_ = lo0073 & new_n5194_;
  assign new_n9311_ = ~new_n9258_ & ~new_n9310_;
  assign new_n9312_ = new_n3936_ & ~new_n9311_;
  assign new_n9313_ = new_n3625_ & new_n9258_;
  assign new_n9314_ = ~new_n9312_ & ~new_n9313_;
  assign new_n9315_ = lo0073 & new_n5608_;
  assign new_n9316_ = ~new_n5184_ & new_n9315_;
  assign new_n9317_ = lo0073 & new_n3706_;
  assign new_n9318_ = ~new_n9309_ & new_n9314_;
  assign new_n9319_ = ~new_n9316_ & new_n9318_;
  assign new_n9320_ = ~new_n9317_ & new_n9319_;
  assign new_n9321_ = new_n5133_ & new_n9308_;
  assign new_n9322_ = new_n9320_ & ~new_n9321_;
  assign new_n9323_ = lo0073 & new_n5505_;
  assign new_n9324_ = new_n9266_ & new_n9307_;
  assign new_n9325_ = new_n9322_ & new_n9324_;
  assign new_n9326_ = ~new_n9323_ & new_n9325_;
  assign new_n9327_ = new_n3804_ & new_n9258_;
  assign new_n9328_ = new_n3834_ & new_n9296_;
  assign new_n9329_ = new_n3678_ & new_n9328_;
  assign new_n9330_ = lo0073 & new_n5112_;
  assign new_n9331_ = new_n3810_ & new_n9276_;
  assign new_n9332_ = ~new_n9327_ & ~new_n9329_;
  assign new_n9333_ = ~new_n9330_ & new_n9332_;
  assign new_n9334_ = ~new_n9331_ & new_n9333_;
  assign new_n9335_ = ~new_n5105_ & new_n9276_;
  assign new_n9336_ = new_n9334_ & ~new_n9335_;
  assign new_n9337_ = new_n3815_ & new_n9257_;
  assign new_n9338_ = new_n4088_ & new_n9258_;
  assign new_n9339_ = ~new_n9337_ & ~new_n9338_;
  assign new_n9340_ = new_n3820_ & new_n9276_;
  assign new_n9341_ = new_n3870_ & new_n9291_;
  assign new_n9342_ = ~new_n9340_ & ~new_n9341_;
  assign new_n9343_ = ~new_n4069_ & new_n9258_;
  assign new_n9344_ = new_n9336_ & new_n9339_;
  assign new_n9345_ = new_n9342_ & new_n9344_;
  assign new_n9346_ = ~new_n9343_ & new_n9345_;
  assign new_n9347_ = new_n4020_ & new_n9258_;
  assign new_n9348_ = ~new_n5096_ & new_n9276_;
  assign new_n9349_ = ~new_n9347_ & ~new_n9348_;
  assign new_n9350_ = ~new_n4096_ & new_n9258_;
  assign new_n9351_ = lo0073 & ~new_n9258_;
  assign new_n9352_ = ~new_n9350_ & ~new_n9351_;
  assign new_n9353_ = new_n5090_ & ~new_n9352_;
  assign new_n9354_ = new_n3746_ & new_n9257_;
  assign new_n9355_ = ~new_n9353_ & ~new_n9354_;
  assign new_n9356_ = lo0073 & new_n5071_;
  assign new_n9357_ = lo0073 & lo0786;
  assign new_n9358_ = lo0073 & new_n5545_;
  assign new_n9359_ = new_n4428_ & new_n4528_;
  assign new_n9360_ = ~new_n5076_ & new_n9296_;
  assign new_n9361_ = ~new_n9359_ & ~new_n9360_;
  assign new_n9362_ = ~new_n9358_ & new_n9361_;
  assign new_n9363_ = new_n4475_ & ~new_n9362_;
  assign new_n9364_ = new_n5082_ & new_n9357_;
  assign new_n9365_ = ~new_n9363_ & ~new_n9364_;
  assign new_n9366_ = ~new_n9356_ & new_n9365_;
  assign new_n9367_ = new_n5070_ & ~new_n9366_;
  assign new_n9368_ = new_n9346_ & new_n9349_;
  assign new_n9369_ = new_n9355_ & new_n9368_;
  assign new_n9370_ = ~new_n9367_ & new_n9369_;
  assign li0073 = ~new_n9326_ | ~new_n9370_;
  assign new_n9372_ = ~lo0024 & lo0074;
  assign new_n9373_ = new_n4050_ & new_n9372_;
  assign new_n9374_ = lo0074 & new_n5562_;
  assign new_n9375_ = lo0074 & ~lo0314;
  assign new_n9376_ = lo0074 & new_n5155_;
  assign new_n9377_ = new_n3777_ & new_n9376_;
  assign new_n9378_ = lo0074 & ~new_n4632_;
  assign new_n9379_ = new_n5565_ & new_n9378_;
  assign new_n9380_ = ~new_n9377_ & ~new_n9379_;
  assign new_n9381_ = ~new_n5460_ & new_n9375_;
  assign new_n9382_ = new_n9380_ & ~new_n9381_;
  assign new_n9383_ = lo0074 & ~lo0841;
  assign new_n9384_ = new_n3763_ & new_n9383_;
  assign new_n9385_ = new_n3780_ & new_n9372_;
  assign new_n9386_ = ~new_n9384_ & ~new_n9385_;
  assign new_n9387_ = new_n3794_ & new_n9375_;
  assign new_n9388_ = new_n9386_ & ~new_n9387_;
  assign new_n9389_ = ~new_n9373_ & ~new_n9374_;
  assign new_n9390_ = new_n9382_ & new_n9389_;
  assign new_n9391_ = new_n9388_ & new_n9390_;
  assign new_n9392_ = new_n4041_ & new_n9372_;
  assign new_n9393_ = new_n9391_ & ~new_n9392_;
  assign new_n9394_ = lo0074 & new_n3678_;
  assign new_n9395_ = new_n3786_ & new_n9372_;
  assign new_n9396_ = new_n5139_ & new_n9394_;
  assign new_n9397_ = ~new_n9395_ & ~new_n9396_;
  assign new_n9398_ = ~lo1044 & new_n9375_;
  assign new_n9399_ = new_n4007_ & new_n9398_;
  assign new_n9400_ = new_n3969_ & new_n9383_;
  assign new_n9401_ = ~new_n9399_ & ~new_n9400_;
  assign new_n9402_ = ~lo0074 & lo0479;
  assign new_n9403_ = ~new_n4053_ & new_n9402_;
  assign new_n9404_ = ~li0583 & ~new_n9403_;
  assign new_n9405_ = lo0074 & li0583;
  assign new_n9406_ = new_n3974_ & ~new_n4135_;
  assign new_n9407_ = ~new_n9404_ & ~new_n9405_;
  assign new_n9408_ = new_n9406_ & ~new_n9407_;
  assign new_n9409_ = new_n4133_ & new_n9372_;
  assign new_n9410_ = ~new_n9408_ & ~new_n9409_;
  assign new_n9411_ = lo0074 & ~new_n5216_;
  assign new_n9412_ = new_n9410_ & ~new_n9411_;
  assign new_n9413_ = new_n3948_ & new_n9372_;
  assign new_n9414_ = new_n9412_ & ~new_n9413_;
  assign new_n9415_ = new_n9393_ & new_n9397_;
  assign new_n9416_ = new_n9401_ & new_n9415_;
  assign new_n9417_ = new_n9414_ & new_n9416_;
  assign new_n9418_ = lo0074 & new_n5505_;
  assign new_n9419_ = lo0074 & new_n5135_;
  assign new_n9420_ = lo0074 & new_n5194_;
  assign new_n9421_ = ~new_n9372_ & ~new_n9420_;
  assign new_n9422_ = new_n3936_ & ~new_n9421_;
  assign new_n9423_ = new_n3625_ & new_n9372_;
  assign new_n9424_ = ~new_n9422_ & ~new_n9423_;
  assign new_n9425_ = lo0074 & new_n3706_;
  assign new_n9426_ = lo0074 & new_n5608_;
  assign new_n9427_ = ~new_n5184_ & new_n9426_;
  assign new_n9428_ = new_n9424_ & ~new_n9425_;
  assign new_n9429_ = ~new_n9427_ & new_n9428_;
  assign new_n9430_ = ~new_n5201_ & new_n9383_;
  assign new_n9431_ = new_n9429_ & ~new_n9430_;
  assign new_n9432_ = ~new_n9418_ & ~new_n9419_;
  assign new_n9433_ = new_n9431_ & new_n9432_;
  assign new_n9434_ = new_n9417_ & new_n9433_;
  assign new_n9435_ = ~new_n5060_ & new_n9375_;
  assign new_n9436_ = new_n3940_ & new_n9372_;
  assign new_n9437_ = ~new_n9435_ & ~new_n9436_;
  assign new_n9438_ = new_n3953_ & new_n9372_;
  assign new_n9439_ = lo0074 & new_n5671_;
  assign new_n9440_ = new_n9437_ & ~new_n9438_;
  assign new_n9441_ = ~new_n9439_ & new_n9440_;
  assign new_n9442_ = ~new_n5105_ & new_n9383_;
  assign new_n9443_ = new_n9441_ & ~new_n9442_;
  assign new_n9444_ = new_n3815_ & new_n9375_;
  assign new_n9445_ = new_n4088_ & new_n9372_;
  assign new_n9446_ = ~new_n9444_ & ~new_n9445_;
  assign new_n9447_ = ~li0683 & ~new_n9402_;
  assign new_n9448_ = lo0841 & new_n9447_;
  assign new_n9449_ = ~new_n9383_ & ~new_n9448_;
  assign new_n9450_ = new_n3810_ & ~new_n9449_;
  assign new_n9451_ = new_n3834_ & new_n9405_;
  assign new_n9452_ = new_n3678_ & new_n9451_;
  assign new_n9453_ = new_n3804_ & new_n9372_;
  assign new_n9454_ = ~new_n9452_ & ~new_n9453_;
  assign new_n9455_ = ~new_n9450_ & new_n9454_;
  assign new_n9456_ = new_n3820_ & new_n9383_;
  assign new_n9457_ = new_n3870_ & new_n9398_;
  assign new_n9458_ = ~new_n9456_ & ~new_n9457_;
  assign new_n9459_ = ~new_n4069_ & new_n9372_;
  assign new_n9460_ = new_n9446_ & new_n9455_;
  assign new_n9461_ = new_n9458_ & new_n9460_;
  assign new_n9462_ = ~new_n9459_ & new_n9461_;
  assign new_n9463_ = new_n4020_ & new_n9372_;
  assign new_n9464_ = ~new_n5096_ & new_n9383_;
  assign new_n9465_ = ~new_n9463_ & ~new_n9464_;
  assign new_n9466_ = lo0074 & new_n5071_;
  assign new_n9467_ = lo0074 & new_n4219_;
  assign new_n9468_ = ~new_n5074_ & new_n9467_;
  assign new_n9469_ = ~new_n5076_ & new_n9405_;
  assign new_n9470_ = ~new_n9468_ & ~new_n9469_;
  assign new_n9471_ = new_n4475_ & ~new_n9470_;
  assign new_n9472_ = lo0074 & new_n5083_;
  assign new_n9473_ = ~new_n9466_ & ~new_n9471_;
  assign new_n9474_ = ~new_n9472_ & new_n9473_;
  assign new_n9475_ = new_n5070_ & ~new_n9474_;
  assign new_n9476_ = ~new_n4096_ & new_n9372_;
  assign new_n9477_ = lo0074 & ~new_n9372_;
  assign new_n9478_ = ~new_n9476_ & ~new_n9477_;
  assign new_n9479_ = new_n5090_ & ~new_n9478_;
  assign new_n9480_ = new_n3746_ & new_n9375_;
  assign new_n9481_ = ~new_n9479_ & ~new_n9480_;
  assign new_n9482_ = new_n9465_ & ~new_n9475_;
  assign new_n9483_ = new_n9481_ & new_n9482_;
  assign new_n9484_ = new_n9462_ & new_n9483_;
  assign new_n9485_ = new_n9434_ & new_n9443_;
  assign li0074 = ~new_n9484_ | ~new_n9485_;
  assign new_n9487_ = lo0075 & ~lo0841;
  assign new_n9488_ = ~lo0024 & lo0075;
  assign new_n9489_ = new_n4020_ & new_n9488_;
  assign new_n9490_ = ~new_n5096_ & new_n9487_;
  assign new_n9491_ = ~new_n9489_ & ~new_n9490_;
  assign new_n9492_ = lo0075 & new_n5071_;
  assign new_n9493_ = lo0075 & new_n4219_;
  assign new_n9494_ = lo0075 & li0583;
  assign new_n9495_ = ~new_n5074_ & new_n9493_;
  assign new_n9496_ = ~new_n5076_ & new_n9494_;
  assign new_n9497_ = ~new_n9495_ & ~new_n9496_;
  assign new_n9498_ = new_n4475_ & ~new_n9497_;
  assign new_n9499_ = lo0075 & new_n5083_;
  assign new_n9500_ = ~new_n9492_ & ~new_n9498_;
  assign new_n9501_ = ~new_n9499_ & new_n9500_;
  assign new_n9502_ = new_n5070_ & ~new_n9501_;
  assign new_n9503_ = ~new_n4096_ & new_n9488_;
  assign new_n9504_ = lo0075 & ~new_n9488_;
  assign new_n9505_ = ~new_n9503_ & ~new_n9504_;
  assign new_n9506_ = lo0075 & ~lo0314;
  assign new_n9507_ = new_n5090_ & ~new_n9505_;
  assign new_n9508_ = new_n3746_ & new_n9506_;
  assign new_n9509_ = ~new_n9507_ & ~new_n9508_;
  assign new_n9510_ = new_n9491_ & ~new_n9502_;
  assign new_n9511_ = new_n9509_ & new_n9510_;
  assign new_n9512_ = lo0075 & new_n5194_;
  assign new_n9513_ = ~new_n9488_ & ~new_n9512_;
  assign new_n9514_ = new_n3936_ & ~new_n9513_;
  assign new_n9515_ = new_n3625_ & new_n9488_;
  assign new_n9516_ = ~new_n9514_ & ~new_n9515_;
  assign new_n9517_ = lo0075 & new_n3706_;
  assign new_n9518_ = lo0075 & new_n5818_;
  assign new_n9519_ = ~new_n5184_ & new_n9518_;
  assign new_n9520_ = new_n9516_ & ~new_n9517_;
  assign new_n9521_ = ~new_n9519_ & new_n9520_;
  assign new_n9522_ = ~new_n5201_ & new_n9487_;
  assign new_n9523_ = new_n9521_ & ~new_n9522_;
  assign new_n9524_ = new_n9511_ & new_n9523_;
  assign new_n9525_ = ~new_n5060_ & new_n9506_;
  assign new_n9526_ = new_n3940_ & new_n9488_;
  assign new_n9527_ = ~new_n9525_ & ~new_n9526_;
  assign new_n9528_ = new_n4050_ & new_n9488_;
  assign new_n9529_ = lo0075 & new_n5562_;
  assign new_n9530_ = lo0075 & new_n5155_;
  assign new_n9531_ = new_n3777_ & new_n9530_;
  assign new_n9532_ = lo0075 & ~new_n4632_;
  assign new_n9533_ = new_n5565_ & new_n9532_;
  assign new_n9534_ = ~new_n9531_ & ~new_n9533_;
  assign new_n9535_ = ~new_n5460_ & new_n9506_;
  assign new_n9536_ = new_n9534_ & ~new_n9535_;
  assign new_n9537_ = new_n3763_ & new_n9487_;
  assign new_n9538_ = new_n3780_ & new_n9488_;
  assign new_n9539_ = ~new_n9537_ & ~new_n9538_;
  assign new_n9540_ = new_n3794_ & new_n9506_;
  assign new_n9541_ = new_n9539_ & ~new_n9540_;
  assign new_n9542_ = ~new_n9528_ & ~new_n9529_;
  assign new_n9543_ = new_n9536_ & new_n9542_;
  assign new_n9544_ = new_n9541_ & new_n9543_;
  assign new_n9545_ = new_n4041_ & new_n9488_;
  assign new_n9546_ = new_n9544_ & ~new_n9545_;
  assign new_n9547_ = lo0075 & ~new_n5216_;
  assign new_n9548_ = new_n4133_ & new_n9488_;
  assign new_n9549_ = ~new_n9547_ & ~new_n9548_;
  assign new_n9550_ = lo0075 & lo0479;
  assign new_n9551_ = new_n5222_ & new_n9550_;
  assign new_n9552_ = ~new_n9494_ & ~new_n9551_;
  assign new_n9553_ = new_n3974_ & ~new_n9552_;
  assign new_n9554_ = new_n3974_ & new_n4135_;
  assign new_n9555_ = new_n9549_ & ~new_n9553_;
  assign new_n9556_ = ~new_n9554_ & new_n9555_;
  assign new_n9557_ = new_n3948_ & new_n9488_;
  assign new_n9558_ = new_n9556_ & ~new_n9557_;
  assign new_n9559_ = lo0075 & new_n3678_;
  assign new_n9560_ = new_n3786_ & new_n9488_;
  assign new_n9561_ = new_n5139_ & new_n9559_;
  assign new_n9562_ = ~new_n9560_ & ~new_n9561_;
  assign new_n9563_ = new_n9527_ & new_n9546_;
  assign new_n9564_ = new_n9558_ & new_n9563_;
  assign new_n9565_ = new_n9562_ & new_n9564_;
  assign new_n9566_ = lo0075 & new_n5135_;
  assign new_n9567_ = ~lo1044 & new_n9506_;
  assign new_n9568_ = new_n4007_ & new_n9567_;
  assign new_n9569_ = new_n3969_ & new_n9487_;
  assign new_n9570_ = ~new_n9568_ & ~new_n9569_;
  assign new_n9571_ = ~new_n9566_ & new_n9570_;
  assign new_n9572_ = lo0075 & new_n5505_;
  assign new_n9573_ = lo0075 & ~lo0993;
  assign new_n9574_ = new_n3927_ & new_n9573_;
  assign new_n9575_ = new_n3953_ & new_n9488_;
  assign new_n9576_ = ~new_n9574_ & ~new_n9575_;
  assign new_n9577_ = new_n9571_ & ~new_n9572_;
  assign new_n9578_ = new_n9576_ & new_n9577_;
  assign new_n9579_ = new_n3834_ & new_n9494_;
  assign new_n9580_ = new_n3678_ & new_n9579_;
  assign new_n9581_ = new_n3804_ & new_n9488_;
  assign new_n9582_ = ~new_n9580_ & ~new_n9581_;
  assign new_n9583_ = ~li0683 & ~new_n9550_;
  assign new_n9584_ = lo0841 & ~new_n9583_;
  assign new_n9585_ = ~new_n9487_ & ~new_n9584_;
  assign new_n9586_ = new_n3810_ & ~new_n9585_;
  assign new_n9587_ = new_n9582_ & ~new_n9586_;
  assign new_n9588_ = ~new_n5105_ & new_n9487_;
  assign new_n9589_ = new_n9587_ & ~new_n9588_;
  assign new_n9590_ = new_n3815_ & new_n9506_;
  assign new_n9591_ = new_n4088_ & new_n9488_;
  assign new_n9592_ = ~new_n9590_ & ~new_n9591_;
  assign new_n9593_ = new_n3820_ & new_n9487_;
  assign new_n9594_ = new_n3870_ & new_n9567_;
  assign new_n9595_ = ~new_n9593_ & ~new_n9594_;
  assign new_n9596_ = ~new_n4069_ & new_n9488_;
  assign new_n9597_ = new_n9589_ & new_n9592_;
  assign new_n9598_ = new_n9595_ & new_n9597_;
  assign new_n9599_ = ~new_n9596_ & new_n9598_;
  assign new_n9600_ = new_n9578_ & new_n9599_;
  assign new_n9601_ = new_n9524_ & new_n9565_;
  assign li0075 = ~new_n9600_ | ~new_n9601_;
  assign new_n9603_ = lo0076 & new_n5505_;
  assign new_n9604_ = ~lo0076 & new_n4647_;
  assign new_n9605_ = new_n3705_ & ~new_n9604_;
  assign new_n9606_ = ~new_n5131_ & new_n9605_;
  assign new_n9607_ = ~new_n5134_ & new_n9606_;
  assign new_n9608_ = lo0076 & ~lo0993;
  assign new_n9609_ = ~lo0024 & lo0076;
  assign new_n9610_ = new_n3927_ & new_n9608_;
  assign new_n9611_ = new_n3953_ & new_n9609_;
  assign new_n9612_ = ~new_n9610_ & ~new_n9611_;
  assign new_n9613_ = lo0076 & ~lo0841;
  assign new_n9614_ = lo0076 & ~lo0314;
  assign new_n9615_ = ~lo1044 & new_n9614_;
  assign new_n9616_ = new_n4007_ & new_n9615_;
  assign new_n9617_ = new_n3969_ & new_n9613_;
  assign new_n9618_ = ~new_n9616_ & ~new_n9617_;
  assign new_n9619_ = ~new_n9603_ & ~new_n9607_;
  assign new_n9620_ = new_n9612_ & new_n9619_;
  assign new_n9621_ = new_n9618_ & new_n9620_;
  assign new_n9622_ = lo0076 & ~new_n5216_;
  assign new_n9623_ = new_n4133_ & new_n9609_;
  assign new_n9624_ = ~new_n9622_ & ~new_n9623_;
  assign new_n9625_ = lo0076 & li0583;
  assign new_n9626_ = new_n3974_ & new_n9625_;
  assign new_n9627_ = ~new_n4135_ & new_n9626_;
  assign new_n9628_ = lo0076 & new_n5225_;
  assign new_n9629_ = new_n9624_ & ~new_n9627_;
  assign new_n9630_ = ~new_n9628_ & new_n9629_;
  assign new_n9631_ = new_n3948_ & new_n9609_;
  assign new_n9632_ = new_n9630_ & ~new_n9631_;
  assign new_n9633_ = lo0076 & new_n3678_;
  assign new_n9634_ = new_n3786_ & new_n9609_;
  assign new_n9635_ = new_n5139_ & new_n9633_;
  assign new_n9636_ = ~new_n9634_ & ~new_n9635_;
  assign new_n9637_ = new_n9632_ & new_n9636_;
  assign new_n9638_ = new_n4050_ & new_n9609_;
  assign new_n9639_ = lo0076 & new_n5562_;
  assign new_n9640_ = lo0076 & new_n5155_;
  assign new_n9641_ = new_n3777_ & new_n9640_;
  assign new_n9642_ = lo0076 & ~new_n4632_;
  assign new_n9643_ = new_n5565_ & new_n9642_;
  assign new_n9644_ = ~new_n9641_ & ~new_n9643_;
  assign new_n9645_ = ~new_n5460_ & new_n9614_;
  assign new_n9646_ = new_n9644_ & ~new_n9645_;
  assign new_n9647_ = new_n3763_ & new_n9613_;
  assign new_n9648_ = new_n3780_ & new_n9609_;
  assign new_n9649_ = ~new_n9647_ & ~new_n9648_;
  assign new_n9650_ = new_n3794_ & new_n9614_;
  assign new_n9651_ = new_n9649_ & ~new_n9650_;
  assign new_n9652_ = ~new_n9638_ & ~new_n9639_;
  assign new_n9653_ = new_n9646_ & new_n9652_;
  assign new_n9654_ = new_n9651_ & new_n9653_;
  assign new_n9655_ = new_n4041_ & new_n9609_;
  assign new_n9656_ = new_n9654_ & ~new_n9655_;
  assign new_n9657_ = lo0076 & new_n5071_;
  assign new_n9658_ = lo0076 & new_n4219_;
  assign new_n9659_ = ~new_n5074_ & new_n9658_;
  assign new_n9660_ = ~new_n5076_ & new_n9625_;
  assign new_n9661_ = ~new_n9659_ & ~new_n9660_;
  assign new_n9662_ = new_n4475_ & ~new_n9661_;
  assign new_n9663_ = lo0076 & new_n5083_;
  assign new_n9664_ = ~new_n9657_ & ~new_n9662_;
  assign new_n9665_ = ~new_n9663_ & new_n9664_;
  assign new_n9666_ = new_n5070_ & ~new_n9665_;
  assign new_n9667_ = ~new_n4096_ & new_n9609_;
  assign new_n9668_ = lo0076 & ~new_n9609_;
  assign new_n9669_ = ~new_n9667_ & ~new_n9668_;
  assign new_n9670_ = new_n5090_ & ~new_n9669_;
  assign new_n9671_ = new_n3746_ & new_n9614_;
  assign new_n9672_ = ~new_n9670_ & ~new_n9671_;
  assign new_n9673_ = new_n9637_ & new_n9656_;
  assign new_n9674_ = ~new_n9666_ & new_n9673_;
  assign new_n9675_ = new_n9672_ & new_n9674_;
  assign new_n9676_ = new_n9621_ & new_n9675_;
  assign new_n9677_ = new_n3804_ & new_n9609_;
  assign new_n9678_ = new_n3834_ & new_n9625_;
  assign new_n9679_ = new_n3678_ & new_n9678_;
  assign new_n9680_ = lo0076 & new_n5112_;
  assign new_n9681_ = new_n3810_ & new_n9613_;
  assign new_n9682_ = ~new_n9677_ & ~new_n9679_;
  assign new_n9683_ = ~new_n9680_ & new_n9682_;
  assign new_n9684_ = ~new_n9681_ & new_n9683_;
  assign new_n9685_ = ~new_n5105_ & new_n9613_;
  assign new_n9686_ = new_n9684_ & ~new_n9685_;
  assign new_n9687_ = lo0076 & new_n5194_;
  assign new_n9688_ = ~new_n9609_ & ~new_n9687_;
  assign new_n9689_ = new_n3936_ & ~new_n9688_;
  assign new_n9690_ = new_n3625_ & new_n9609_;
  assign new_n9691_ = ~new_n9689_ & ~new_n9690_;
  assign new_n9692_ = lo0076 & new_n3706_;
  assign new_n9693_ = lo0076 & new_n5818_;
  assign new_n9694_ = ~new_n5184_ & new_n9693_;
  assign new_n9695_ = new_n9691_ & ~new_n9692_;
  assign new_n9696_ = ~new_n9694_ & new_n9695_;
  assign new_n9697_ = ~new_n5201_ & new_n9613_;
  assign new_n9698_ = new_n9696_ & ~new_n9697_;
  assign new_n9699_ = new_n4020_ & new_n9609_;
  assign new_n9700_ = ~new_n5096_ & new_n9613_;
  assign new_n9701_ = ~new_n9699_ & ~new_n9700_;
  assign new_n9702_ = ~new_n5060_ & new_n9614_;
  assign new_n9703_ = new_n3940_ & new_n9609_;
  assign new_n9704_ = ~new_n9702_ & ~new_n9703_;
  assign new_n9705_ = new_n9701_ & new_n9704_;
  assign new_n9706_ = new_n3815_ & new_n9614_;
  assign new_n9707_ = new_n4088_ & new_n9609_;
  assign new_n9708_ = ~new_n9706_ & ~new_n9707_;
  assign new_n9709_ = ~new_n4069_ & new_n9609_;
  assign new_n9710_ = new_n3820_ & new_n9613_;
  assign new_n9711_ = new_n3870_ & new_n9615_;
  assign new_n9712_ = ~new_n9710_ & ~new_n9711_;
  assign new_n9713_ = new_n9708_ & ~new_n9709_;
  assign new_n9714_ = new_n9712_ & new_n9713_;
  assign new_n9715_ = new_n9705_ & new_n9714_;
  assign new_n9716_ = new_n9686_ & new_n9698_;
  assign new_n9717_ = new_n9715_ & new_n9716_;
  assign li0076 = ~new_n9676_ | ~new_n9717_;
  assign new_n9719_ = lo0077 & ~lo0841;
  assign new_n9720_ = ~lo0024 & lo0077;
  assign new_n9721_ = new_n4020_ & new_n9720_;
  assign new_n9722_ = ~new_n5096_ & new_n9719_;
  assign new_n9723_ = ~new_n9721_ & ~new_n9722_;
  assign new_n9724_ = lo0077 & new_n5071_;
  assign new_n9725_ = lo0077 & li0583;
  assign new_n9726_ = lo0077 & new_n4219_;
  assign new_n9727_ = ~new_n5076_ & new_n9725_;
  assign new_n9728_ = ~new_n5074_ & new_n9726_;
  assign new_n9729_ = ~new_n9727_ & ~new_n9728_;
  assign new_n9730_ = new_n4475_ & ~new_n9729_;
  assign new_n9731_ = lo0077 & new_n5083_;
  assign new_n9732_ = ~new_n9724_ & ~new_n9730_;
  assign new_n9733_ = ~new_n9731_ & new_n9732_;
  assign new_n9734_ = new_n5070_ & ~new_n9733_;
  assign new_n9735_ = ~new_n4096_ & new_n9720_;
  assign new_n9736_ = lo0077 & ~new_n9720_;
  assign new_n9737_ = ~new_n9735_ & ~new_n9736_;
  assign new_n9738_ = lo0077 & ~lo0314;
  assign new_n9739_ = new_n5090_ & ~new_n9737_;
  assign new_n9740_ = new_n3746_ & new_n9738_;
  assign new_n9741_ = ~new_n9739_ & ~new_n9740_;
  assign new_n9742_ = new_n9723_ & ~new_n9734_;
  assign new_n9743_ = new_n9741_ & new_n9742_;
  assign new_n9744_ = lo0077 & ~lo0993;
  assign new_n9745_ = new_n3927_ & new_n9744_;
  assign new_n9746_ = new_n3953_ & new_n9720_;
  assign new_n9747_ = ~new_n9745_ & ~new_n9746_;
  assign new_n9748_ = new_n3763_ & new_n9719_;
  assign new_n9749_ = new_n3780_ & new_n9720_;
  assign new_n9750_ = ~new_n9748_ & ~new_n9749_;
  assign new_n9751_ = new_n3794_ & new_n9738_;
  assign new_n9752_ = new_n9750_ & ~new_n9751_;
  assign new_n9753_ = ~new_n5460_ & new_n9738_;
  assign new_n9754_ = lo0077 & ~new_n4632_;
  assign new_n9755_ = new_n5565_ & new_n9754_;
  assign new_n9756_ = lo0077 & new_n6643_;
  assign new_n9757_ = new_n9752_ & ~new_n9753_;
  assign new_n9758_ = ~new_n9755_ & new_n9757_;
  assign new_n9759_ = ~new_n9756_ & new_n9758_;
  assign new_n9760_ = ~new_n3799_ & new_n9759_;
  assign new_n9761_ = lo0077 & new_n5562_;
  assign new_n9762_ = new_n4050_ & new_n9720_;
  assign new_n9763_ = ~new_n9761_ & ~new_n9762_;
  assign new_n9764_ = new_n4041_ & new_n9720_;
  assign new_n9765_ = new_n9763_ & ~new_n9764_;
  assign new_n9766_ = lo0077 & new_n5140_;
  assign new_n9767_ = new_n3786_ & new_n9720_;
  assign new_n9768_ = new_n9760_ & new_n9765_;
  assign new_n9769_ = ~new_n9766_ & new_n9768_;
  assign new_n9770_ = ~new_n9767_ & new_n9769_;
  assign new_n9771_ = new_n3948_ & new_n9720_;
  assign new_n9772_ = new_n9770_ & ~new_n9771_;
  assign new_n9773_ = ~lo1044 & new_n9738_;
  assign new_n9774_ = new_n4007_ & new_n9773_;
  assign new_n9775_ = new_n3969_ & new_n9719_;
  assign new_n9776_ = ~new_n9774_ & ~new_n9775_;
  assign new_n9777_ = lo0077 & ~new_n5216_;
  assign new_n9778_ = new_n4133_ & new_n9720_;
  assign new_n9779_ = ~new_n9777_ & ~new_n9778_;
  assign new_n9780_ = ~new_n4135_ & new_n9725_;
  assign new_n9781_ = new_n3974_ & new_n9780_;
  assign new_n9782_ = lo0077 & ~new_n4135_;
  assign new_n9783_ = new_n5224_ & new_n9782_;
  assign new_n9784_ = ~new_n9781_ & ~new_n9783_;
  assign new_n9785_ = new_n9779_ & new_n9784_;
  assign new_n9786_ = new_n9747_ & new_n9772_;
  assign new_n9787_ = new_n9776_ & new_n9786_;
  assign new_n9788_ = new_n9785_ & new_n9787_;
  assign new_n9789_ = new_n3804_ & new_n9720_;
  assign new_n9790_ = new_n3834_ & new_n9725_;
  assign new_n9791_ = new_n3678_ & new_n9790_;
  assign new_n9792_ = lo0077 & new_n5112_;
  assign new_n9793_ = new_n3810_ & new_n9719_;
  assign new_n9794_ = ~new_n9789_ & ~new_n9791_;
  assign new_n9795_ = ~new_n9792_ & new_n9794_;
  assign new_n9796_ = ~new_n9793_ & new_n9795_;
  assign new_n9797_ = ~new_n5105_ & new_n9719_;
  assign new_n9798_ = new_n9796_ & ~new_n9797_;
  assign new_n9799_ = new_n3815_ & new_n9738_;
  assign new_n9800_ = new_n4088_ & new_n9720_;
  assign new_n9801_ = ~new_n9799_ & ~new_n9800_;
  assign new_n9802_ = new_n3820_ & new_n9719_;
  assign new_n9803_ = new_n3870_ & new_n9773_;
  assign new_n9804_ = ~new_n9802_ & ~new_n9803_;
  assign new_n9805_ = ~new_n4069_ & new_n9720_;
  assign new_n9806_ = new_n9798_ & new_n9801_;
  assign new_n9807_ = new_n9804_ & new_n9806_;
  assign new_n9808_ = ~new_n9805_ & new_n9807_;
  assign new_n9809_ = lo0077 & new_n5135_;
  assign new_n9810_ = new_n3940_ & new_n9720_;
  assign new_n9811_ = ~new_n9809_ & ~new_n9810_;
  assign new_n9812_ = ~new_n5060_ & new_n9738_;
  assign new_n9813_ = new_n9811_ & ~new_n9812_;
  assign new_n9814_ = lo0077 & new_n5505_;
  assign new_n9815_ = lo0077 & new_n5194_;
  assign new_n9816_ = ~new_n9720_ & ~new_n9815_;
  assign new_n9817_ = new_n3936_ & ~new_n9816_;
  assign new_n9818_ = new_n3625_ & new_n9720_;
  assign new_n9819_ = ~new_n9817_ & ~new_n9818_;
  assign new_n9820_ = lo0077 & new_n3706_;
  assign new_n9821_ = lo0077 & new_n5708_;
  assign new_n9822_ = new_n9819_ & ~new_n9820_;
  assign new_n9823_ = ~new_n9821_ & new_n9822_;
  assign new_n9824_ = ~new_n5201_ & new_n9719_;
  assign new_n9825_ = new_n9823_ & ~new_n9824_;
  assign new_n9826_ = new_n9813_ & ~new_n9814_;
  assign new_n9827_ = new_n9825_ & new_n9826_;
  assign new_n9828_ = new_n9743_ & new_n9788_;
  assign new_n9829_ = new_n9808_ & new_n9828_;
  assign li0077 = ~new_n9827_ | ~new_n9829_;
  assign new_n9831_ = lo0232 & ~lo0468;
  assign li0078 = lo0119 & new_n9831_;
  assign new_n9833_ = ~lo0074 & ~new_n4523_;
  assign new_n9834_ = new_n5259_ & new_n9833_;
  assign new_n9835_ = lo0187 & ~new_n3522_;
  assign new_n9836_ = lo0147 & ~lo0187;
  assign new_n9837_ = ~new_n9835_ & ~new_n9836_;
  assign new_n9838_ = new_n4543_ & new_n9837_;
  assign new_n9839_ = ~lo0040 & new_n5268_;
  assign new_n9840_ = ~lo0079 & new_n5325_;
  assign new_n9841_ = lo0079 & ~new_n5325_;
  assign new_n9842_ = ~new_n9840_ & ~new_n9841_;
  assign new_n9843_ = new_n5276_ & ~new_n9842_;
  assign new_n9844_ = lo0079 & ~new_n5276_;
  assign new_n9845_ = ~new_n9843_ & ~new_n9844_;
  assign new_n9846_ = new_n3579_ & new_n9845_;
  assign new_n9847_ = ~new_n5268_ & ~new_n9838_;
  assign new_n9848_ = new_n9839_ & ~new_n9846_;
  assign new_n9849_ = ~new_n9847_ & ~new_n9848_;
  assign new_n9850_ = lo0184 & ~new_n3522_;
  assign new_n9851_ = lo0163 & ~lo0184;
  assign new_n9852_ = ~new_n9850_ & ~new_n9851_;
  assign new_n9853_ = new_n4543_ & new_n9852_;
  assign new_n9854_ = ~new_n5259_ & ~new_n9853_;
  assign new_n9855_ = ~new_n4553_ & new_n5289_;
  assign new_n9856_ = ~new_n9854_ & ~new_n9855_;
  assign new_n9857_ = new_n9834_ & ~new_n9849_;
  assign new_n9858_ = new_n9856_ & ~new_n9857_;
  assign new_n9859_ = ~new_n5292_ & ~new_n5301_;
  assign new_n9860_ = new_n4543_ & ~new_n9859_;
  assign new_n9861_ = ~new_n5354_ & ~new_n9860_;
  assign new_n9862_ = ~new_n5353_ & ~new_n9861_;
  assign new_n9863_ = ~new_n9853_ & new_n9862_;
  assign new_n9864_ = new_n9853_ & ~new_n9862_;
  assign new_n9865_ = ~new_n9863_ & ~new_n9864_;
  assign new_n9866_ = ~new_n5297_ & ~new_n9858_;
  assign new_n9867_ = new_n9858_ & ~new_n9865_;
  assign new_n9868_ = ~new_n9866_ & ~new_n9867_;
  assign new_n9869_ = ~new_n5252_ & ~new_n6037_;
  assign new_n9870_ = new_n5252_ & ~new_n9868_;
  assign new_n9871_ = ~new_n9869_ & ~new_n9870_;
  assign new_n9872_ = new_n5313_ & new_n9871_;
  assign new_n9873_ = new_n3525_ & ~new_n5313_;
  assign new_n9874_ = ~new_n9872_ & ~new_n9873_;
  assign new_n9875_ = new_n5245_ & ~new_n5317_;
  assign new_n9876_ = lo0179 & ~new_n3522_;
  assign new_n9877_ = lo0156 & ~lo0179;
  assign new_n9878_ = ~new_n9876_ & ~new_n9877_;
  assign new_n9879_ = ~new_n5245_ & new_n9878_;
  assign new_n9880_ = ~new_n9874_ & new_n9875_;
  assign new_n9881_ = ~new_n9879_ & ~new_n9880_;
  assign li0079 = new_n5321_ | new_n9881_;
  assign new_n9883_ = ~lo0080 & new_n5051_;
  assign li0080 = ~new_n5049_ & new_n9883_;
  assign new_n9885_ = lo0081 & ~lo0841;
  assign new_n9886_ = ~lo0024 & lo0081;
  assign new_n9887_ = new_n3804_ & new_n9886_;
  assign new_n9888_ = lo0081 & li0583;
  assign new_n9889_ = new_n3834_ & new_n9888_;
  assign new_n9890_ = new_n3678_ & new_n9889_;
  assign new_n9891_ = lo0081 & new_n5112_;
  assign new_n9892_ = new_n3810_ & new_n9885_;
  assign new_n9893_ = ~new_n9887_ & ~new_n9890_;
  assign new_n9894_ = ~new_n9891_ & new_n9893_;
  assign new_n9895_ = ~new_n9892_ & new_n9894_;
  assign new_n9896_ = ~new_n4069_ & new_n9886_;
  assign new_n9897_ = new_n9895_ & ~new_n9896_;
  assign new_n9898_ = lo0081 & ~lo0314;
  assign new_n9899_ = ~lo1044 & new_n9898_;
  assign new_n9900_ = new_n3820_ & new_n9885_;
  assign new_n9901_ = new_n3870_ & new_n9899_;
  assign new_n9902_ = ~new_n9900_ & ~new_n9901_;
  assign new_n9903_ = new_n9897_ & new_n9902_;
  assign new_n9904_ = ~new_n5105_ & new_n9885_;
  assign new_n9905_ = new_n9903_ & ~new_n9904_;
  assign new_n9906_ = lo0081 & ~new_n5216_;
  assign new_n9907_ = new_n4133_ & new_n9886_;
  assign new_n9908_ = ~new_n9906_ & ~new_n9907_;
  assign new_n9909_ = new_n3974_ & new_n9888_;
  assign new_n9910_ = ~new_n4135_ & new_n9909_;
  assign new_n9911_ = lo0081 & new_n5225_;
  assign new_n9912_ = new_n9908_ & ~new_n9910_;
  assign new_n9913_ = ~new_n9911_ & new_n9912_;
  assign new_n9914_ = new_n3948_ & new_n9886_;
  assign new_n9915_ = new_n9913_ & ~new_n9914_;
  assign new_n9916_ = lo0081 & new_n5671_;
  assign new_n9917_ = lo0081 & new_n3678_;
  assign new_n9918_ = new_n3786_ & new_n9886_;
  assign new_n9919_ = new_n5139_ & new_n9917_;
  assign new_n9920_ = ~new_n9918_ & ~new_n9919_;
  assign new_n9921_ = new_n9905_ & new_n9915_;
  assign new_n9922_ = ~new_n9916_ & new_n9921_;
  assign new_n9923_ = new_n9920_ & new_n9922_;
  assign new_n9924_ = new_n4050_ & new_n9886_;
  assign new_n9925_ = lo0081 & new_n5562_;
  assign new_n9926_ = lo0081 & new_n5155_;
  assign new_n9927_ = new_n3777_ & new_n9926_;
  assign new_n9928_ = lo0081 & ~new_n4632_;
  assign new_n9929_ = new_n5565_ & new_n9928_;
  assign new_n9930_ = ~new_n9927_ & ~new_n9929_;
  assign new_n9931_ = ~new_n5460_ & new_n9898_;
  assign new_n9932_ = new_n9930_ & ~new_n9931_;
  assign new_n9933_ = new_n3763_ & new_n9885_;
  assign new_n9934_ = new_n3780_ & new_n9886_;
  assign new_n9935_ = ~new_n9933_ & ~new_n9934_;
  assign new_n9936_ = new_n3794_ & new_n9898_;
  assign new_n9937_ = new_n9935_ & ~new_n9936_;
  assign new_n9938_ = ~new_n9924_ & ~new_n9925_;
  assign new_n9939_ = new_n9932_ & new_n9938_;
  assign new_n9940_ = new_n9937_ & new_n9939_;
  assign new_n9941_ = new_n4041_ & new_n9886_;
  assign new_n9942_ = new_n9940_ & ~new_n9941_;
  assign new_n9943_ = lo0081 & new_n5194_;
  assign new_n9944_ = ~new_n9886_ & ~new_n9943_;
  assign new_n9945_ = new_n3936_ & ~new_n9944_;
  assign new_n9946_ = new_n3625_ & new_n9886_;
  assign new_n9947_ = ~new_n9945_ & ~new_n9946_;
  assign new_n9948_ = lo0081 & new_n3706_;
  assign new_n9949_ = lo0081 & new_n5818_;
  assign new_n9950_ = ~new_n5184_ & new_n9949_;
  assign new_n9951_ = new_n9947_ & ~new_n9948_;
  assign new_n9952_ = ~new_n9950_ & new_n9951_;
  assign new_n9953_ = ~new_n5096_ & new_n9885_;
  assign new_n9954_ = new_n4020_ & new_n9886_;
  assign new_n9955_ = ~new_n9953_ & ~new_n9954_;
  assign new_n9956_ = lo0081 & new_n5071_;
  assign new_n9957_ = lo0081 & lo0786;
  assign new_n9958_ = ~new_n5076_ & new_n9888_;
  assign new_n9959_ = lo0081 & new_n5545_;
  assign new_n9960_ = ~new_n9958_ & ~new_n9959_;
  assign new_n9961_ = new_n4475_ & ~new_n9960_;
  assign new_n9962_ = new_n5082_ & new_n9957_;
  assign new_n9963_ = ~new_n9961_ & ~new_n9962_;
  assign new_n9964_ = ~new_n9956_ & new_n9963_;
  assign new_n9965_ = new_n5070_ & ~new_n9964_;
  assign new_n9966_ = new_n3746_ & new_n9898_;
  assign new_n9967_ = ~new_n4096_ & new_n9886_;
  assign new_n9968_ = lo0081 & ~new_n9886_;
  assign new_n9969_ = ~new_n9967_ & ~new_n9968_;
  assign new_n9970_ = new_n5090_ & ~new_n9969_;
  assign new_n9971_ = ~new_n9966_ & ~new_n9970_;
  assign new_n9972_ = ~new_n9965_ & new_n9971_;
  assign new_n9973_ = new_n9955_ & new_n9972_;
  assign new_n9974_ = new_n9952_ & new_n9973_;
  assign new_n9975_ = lo0081 & new_n4001_;
  assign new_n9976_ = ~new_n5060_ & new_n9898_;
  assign new_n9977_ = new_n3940_ & new_n9886_;
  assign new_n9978_ = ~new_n9976_ & ~new_n9977_;
  assign new_n9979_ = new_n3953_ & new_n9886_;
  assign new_n9980_ = new_n3815_ & new_n9898_;
  assign new_n9981_ = new_n4088_ & new_n9886_;
  assign new_n9982_ = ~new_n9980_ & ~new_n9981_;
  assign new_n9983_ = new_n9978_ & ~new_n9979_;
  assign new_n9984_ = new_n9982_ & new_n9983_;
  assign new_n9985_ = ~new_n3828_ & new_n9984_;
  assign new_n9986_ = lo0081 & new_n5133_;
  assign new_n9987_ = ~new_n5134_ & new_n9986_;
  assign new_n9988_ = new_n4007_ & new_n9899_;
  assign new_n9989_ = new_n3969_ & new_n9885_;
  assign new_n9990_ = ~new_n9988_ & ~new_n9989_;
  assign new_n9991_ = ~new_n5201_ & new_n9885_;
  assign new_n9992_ = new_n9985_ & ~new_n9987_;
  assign new_n9993_ = new_n9990_ & new_n9992_;
  assign new_n9994_ = ~new_n9991_ & new_n9993_;
  assign new_n9995_ = new_n5230_ & new_n9975_;
  assign new_n9996_ = new_n9994_ & ~new_n9995_;
  assign new_n9997_ = new_n9923_ & new_n9942_;
  assign new_n9998_ = new_n9974_ & new_n9997_;
  assign li0081 = ~new_n9996_ | ~new_n9998_;
  assign new_n10000_ = lo0082 & ~lo0841;
  assign new_n10001_ = lo0082 & new_n5505_;
  assign new_n10002_ = ~new_n5201_ & new_n10000_;
  assign new_n10003_ = ~new_n10001_ & ~new_n10002_;
  assign new_n10004_ = lo0082 & new_n5135_;
  assign new_n10005_ = ~lo0024 & lo0082;
  assign new_n10006_ = new_n3780_ & new_n10005_;
  assign new_n10007_ = new_n3763_ & new_n10000_;
  assign new_n10008_ = ~new_n10006_ & ~new_n10007_;
  assign new_n10009_ = new_n10003_ & ~new_n10004_;
  assign new_n10010_ = new_n10008_ & new_n10009_;
  assign new_n10011_ = new_n3804_ & new_n10005_;
  assign new_n10012_ = lo0082 & li0583;
  assign new_n10013_ = new_n3834_ & new_n10012_;
  assign new_n10014_ = new_n3678_ & new_n10013_;
  assign new_n10015_ = lo0082 & new_n5112_;
  assign new_n10016_ = new_n3810_ & new_n10000_;
  assign new_n10017_ = ~new_n10011_ & ~new_n10014_;
  assign new_n10018_ = ~new_n10015_ & new_n10017_;
  assign new_n10019_ = ~new_n10016_ & new_n10018_;
  assign new_n10020_ = ~new_n4069_ & new_n10005_;
  assign new_n10021_ = new_n10019_ & ~new_n10020_;
  assign new_n10022_ = lo0082 & ~lo0314;
  assign new_n10023_ = ~lo1044 & new_n10022_;
  assign new_n10024_ = new_n3820_ & new_n10000_;
  assign new_n10025_ = new_n3870_ & new_n10023_;
  assign new_n10026_ = ~new_n10024_ & ~new_n10025_;
  assign new_n10027_ = new_n10021_ & new_n10026_;
  assign new_n10028_ = ~new_n5105_ & new_n10000_;
  assign new_n10029_ = new_n10027_ & ~new_n10028_;
  assign new_n10030_ = lo0082 & new_n5194_;
  assign new_n10031_ = ~new_n10005_ & ~new_n10030_;
  assign new_n10032_ = new_n3936_ & ~new_n10031_;
  assign new_n10033_ = new_n3625_ & new_n10005_;
  assign new_n10034_ = ~new_n10032_ & ~new_n10033_;
  assign new_n10035_ = lo0082 & new_n3706_;
  assign new_n10036_ = lo0082 & new_n5818_;
  assign new_n10037_ = ~new_n5184_ & new_n10036_;
  assign new_n10038_ = new_n10034_ & ~new_n10035_;
  assign new_n10039_ = ~new_n10037_ & new_n10038_;
  assign new_n10040_ = ~new_n5096_ & new_n10000_;
  assign new_n10041_ = new_n4020_ & new_n10005_;
  assign new_n10042_ = ~new_n10040_ & ~new_n10041_;
  assign new_n10043_ = lo0082 & new_n5071_;
  assign new_n10044_ = lo0082 & lo0786;
  assign new_n10045_ = ~new_n5076_ & new_n10012_;
  assign new_n10046_ = lo0082 & new_n5545_;
  assign new_n10047_ = ~new_n10045_ & ~new_n10046_;
  assign new_n10048_ = new_n4475_ & ~new_n10047_;
  assign new_n10049_ = new_n5082_ & new_n10044_;
  assign new_n10050_ = ~new_n10048_ & ~new_n10049_;
  assign new_n10051_ = ~new_n10043_ & new_n10050_;
  assign new_n10052_ = new_n5070_ & ~new_n10051_;
  assign new_n10053_ = new_n3746_ & new_n10022_;
  assign new_n10054_ = ~new_n4096_ & new_n10005_;
  assign new_n10055_ = lo0082 & ~new_n10005_;
  assign new_n10056_ = ~new_n10054_ & ~new_n10055_;
  assign new_n10057_ = new_n5090_ & ~new_n10056_;
  assign new_n10058_ = ~new_n10053_ & ~new_n10057_;
  assign new_n10059_ = ~new_n10052_ & new_n10058_;
  assign new_n10060_ = new_n10042_ & new_n10059_;
  assign new_n10061_ = new_n10029_ & new_n10039_;
  assign new_n10062_ = new_n10060_ & new_n10061_;
  assign new_n10063_ = new_n10010_ & new_n10062_;
  assign new_n10064_ = new_n4050_ & new_n10005_;
  assign new_n10065_ = lo0082 & new_n3678_;
  assign new_n10066_ = new_n5139_ & new_n10065_;
  assign new_n10067_ = new_n3948_ & new_n10005_;
  assign new_n10068_ = ~new_n10066_ & ~new_n10067_;
  assign new_n10069_ = new_n3969_ & new_n10000_;
  assign new_n10070_ = new_n10068_ & ~new_n10069_;
  assign new_n10071_ = new_n4007_ & new_n10023_;
  assign new_n10072_ = lo0082 & new_n5562_;
  assign new_n10073_ = ~new_n10064_ & new_n10070_;
  assign new_n10074_ = ~new_n10071_ & new_n10073_;
  assign new_n10075_ = ~new_n10072_ & new_n10074_;
  assign new_n10076_ = new_n3786_ & new_n10005_;
  assign new_n10077_ = lo0082 & ~new_n5216_;
  assign new_n10078_ = new_n4133_ & new_n10005_;
  assign new_n10079_ = ~new_n10077_ & ~new_n10078_;
  assign new_n10080_ = new_n3974_ & new_n10012_;
  assign new_n10081_ = ~new_n4135_ & new_n10080_;
  assign new_n10082_ = lo0082 & new_n5225_;
  assign new_n10083_ = new_n10079_ & ~new_n10081_;
  assign new_n10084_ = ~new_n10082_ & new_n10083_;
  assign new_n10085_ = ~new_n10076_ & new_n10084_;
  assign new_n10086_ = new_n10075_ & new_n10085_;
  assign new_n10087_ = ~new_n5060_ & new_n10022_;
  assign new_n10088_ = new_n3940_ & new_n10005_;
  assign new_n10089_ = ~new_n10087_ & ~new_n10088_;
  assign new_n10090_ = new_n3815_ & new_n10022_;
  assign new_n10091_ = new_n4088_ & new_n10005_;
  assign new_n10092_ = ~new_n10090_ & ~new_n10091_;
  assign new_n10093_ = new_n3953_ & new_n10005_;
  assign new_n10094_ = new_n10089_ & new_n10092_;
  assign new_n10095_ = ~new_n10093_ & new_n10094_;
  assign new_n10096_ = ~new_n3846_ & new_n10095_;
  assign new_n10097_ = ~lo0082 & ~lo0314;
  assign new_n10098_ = new_n3794_ & ~new_n10097_;
  assign new_n10099_ = new_n3903_ & new_n10022_;
  assign new_n10100_ = ~new_n10098_ & ~new_n10099_;
  assign new_n10101_ = lo0082 & new_n6643_;
  assign new_n10102_ = lo0082 & ~new_n4632_;
  assign new_n10103_ = new_n5565_ & new_n10102_;
  assign new_n10104_ = new_n10100_ & ~new_n10101_;
  assign new_n10105_ = ~new_n10103_ & new_n10104_;
  assign new_n10106_ = new_n3914_ & new_n10022_;
  assign new_n10107_ = new_n10105_ & ~new_n10106_;
  assign new_n10108_ = lo0082 & new_n5671_;
  assign new_n10109_ = new_n4041_ & new_n10005_;
  assign new_n10110_ = new_n10107_ & ~new_n10108_;
  assign new_n10111_ = ~new_n10109_ & new_n10110_;
  assign new_n10112_ = new_n10096_ & new_n10111_;
  assign new_n10113_ = new_n10086_ & new_n10112_;
  assign li0082 = ~new_n10063_ | ~new_n10113_;
  assign new_n10115_ = lo0083 & ~new_n5134_;
  assign new_n10116_ = lo0083 & new_n5230_;
  assign new_n10117_ = new_n4001_ & new_n10116_;
  assign new_n10118_ = new_n5133_ & new_n10115_;
  assign new_n10119_ = ~new_n10117_ & ~new_n10118_;
  assign new_n10120_ = lo0083 & new_n5818_;
  assign new_n10121_ = ~new_n5184_ & new_n10120_;
  assign new_n10122_ = ~lo0024 & lo0083;
  assign new_n10123_ = lo0083 & new_n5194_;
  assign new_n10124_ = ~new_n10122_ & ~new_n10123_;
  assign new_n10125_ = new_n3936_ & ~new_n10124_;
  assign new_n10126_ = new_n3625_ & new_n10122_;
  assign new_n10127_ = ~new_n10125_ & ~new_n10126_;
  assign new_n10128_ = lo0083 & ~lo0841;
  assign new_n10129_ = ~new_n5201_ & new_n10128_;
  assign new_n10130_ = lo0083 & new_n3706_;
  assign new_n10131_ = ~new_n10121_ & new_n10127_;
  assign new_n10132_ = ~new_n10129_ & new_n10131_;
  assign new_n10133_ = ~new_n10130_ & new_n10132_;
  assign new_n10134_ = lo0083 & ~lo0314;
  assign new_n10135_ = ~new_n5060_ & new_n10134_;
  assign new_n10136_ = new_n3940_ & new_n10122_;
  assign new_n10137_ = ~new_n10135_ & ~new_n10136_;
  assign new_n10138_ = lo0083 & ~lo0993;
  assign new_n10139_ = new_n3927_ & new_n10138_;
  assign new_n10140_ = new_n3953_ & new_n10122_;
  assign new_n10141_ = ~new_n10139_ & ~new_n10140_;
  assign new_n10142_ = new_n10137_ & new_n10141_;
  assign new_n10143_ = ~lo1044 & new_n10134_;
  assign new_n10144_ = new_n4007_ & new_n10143_;
  assign new_n10145_ = new_n3969_ & new_n10128_;
  assign new_n10146_ = ~new_n10144_ & ~new_n10145_;
  assign new_n10147_ = new_n3948_ & new_n10122_;
  assign new_n10148_ = lo0083 & li0583;
  assign new_n10149_ = new_n3974_ & new_n10148_;
  assign new_n10150_ = ~new_n4135_ & new_n10149_;
  assign new_n10151_ = lo0083 & new_n5225_;
  assign new_n10152_ = ~new_n10150_ & ~new_n10151_;
  assign new_n10153_ = lo0083 & ~new_n5216_;
  assign new_n10154_ = new_n4133_ & new_n10122_;
  assign new_n10155_ = ~new_n10153_ & ~new_n10154_;
  assign new_n10156_ = new_n10146_ & ~new_n10147_;
  assign new_n10157_ = new_n10152_ & new_n10156_;
  assign new_n10158_ = new_n10155_ & new_n10157_;
  assign new_n10159_ = new_n10142_ & new_n10158_;
  assign new_n10160_ = lo0083 & new_n5155_;
  assign new_n10161_ = new_n3777_ & new_n10160_;
  assign new_n10162_ = lo0083 & ~new_n4632_;
  assign new_n10163_ = new_n5565_ & new_n10162_;
  assign new_n10164_ = ~new_n10161_ & ~new_n10163_;
  assign new_n10165_ = ~new_n5460_ & new_n10134_;
  assign new_n10166_ = new_n10164_ & ~new_n10165_;
  assign new_n10167_ = lo0083 & new_n5562_;
  assign new_n10168_ = new_n4050_ & new_n10122_;
  assign new_n10169_ = new_n3763_ & new_n10128_;
  assign new_n10170_ = new_n3780_ & new_n10122_;
  assign new_n10171_ = ~new_n10169_ & ~new_n10170_;
  assign new_n10172_ = new_n3794_ & new_n10134_;
  assign new_n10173_ = new_n10171_ & ~new_n10172_;
  assign new_n10174_ = new_n10166_ & ~new_n10167_;
  assign new_n10175_ = ~new_n10168_ & new_n10174_;
  assign new_n10176_ = new_n10173_ & new_n10175_;
  assign new_n10177_ = new_n4041_ & new_n10122_;
  assign new_n10178_ = new_n10176_ & ~new_n10177_;
  assign new_n10179_ = new_n3786_ & new_n10122_;
  assign new_n10180_ = lo0083 & new_n5140_;
  assign new_n10181_ = new_n10178_ & ~new_n10179_;
  assign new_n10182_ = ~new_n10180_ & new_n10181_;
  assign new_n10183_ = new_n10119_ & new_n10133_;
  assign new_n10184_ = new_n10159_ & new_n10183_;
  assign new_n10185_ = new_n10182_ & new_n10184_;
  assign new_n10186_ = ~new_n5096_ & new_n10128_;
  assign new_n10187_ = new_n4020_ & new_n10122_;
  assign new_n10188_ = ~new_n10186_ & ~new_n10187_;
  assign new_n10189_ = lo0083 & new_n5071_;
  assign new_n10190_ = lo0083 & lo0786;
  assign new_n10191_ = ~new_n5076_ & new_n10148_;
  assign new_n10192_ = lo0083 & new_n5545_;
  assign new_n10193_ = ~new_n10191_ & ~new_n10192_;
  assign new_n10194_ = new_n4475_ & ~new_n10193_;
  assign new_n10195_ = new_n5082_ & new_n10190_;
  assign new_n10196_ = ~new_n10194_ & ~new_n10195_;
  assign new_n10197_ = ~new_n10189_ & new_n10196_;
  assign new_n10198_ = new_n5070_ & ~new_n10197_;
  assign new_n10199_ = new_n3746_ & new_n10134_;
  assign new_n10200_ = ~new_n4096_ & new_n10122_;
  assign new_n10201_ = lo0083 & ~new_n10122_;
  assign new_n10202_ = ~new_n10200_ & ~new_n10201_;
  assign new_n10203_ = new_n5090_ & ~new_n10202_;
  assign new_n10204_ = ~new_n10199_ & ~new_n10203_;
  assign new_n10205_ = ~new_n10198_ & new_n10204_;
  assign new_n10206_ = new_n10188_ & new_n10205_;
  assign new_n10207_ = new_n3804_ & new_n10122_;
  assign new_n10208_ = new_n3834_ & new_n10148_;
  assign new_n10209_ = new_n3678_ & new_n10208_;
  assign new_n10210_ = lo0083 & new_n5112_;
  assign new_n10211_ = new_n3810_ & new_n10128_;
  assign new_n10212_ = ~new_n10207_ & ~new_n10209_;
  assign new_n10213_ = ~new_n10210_ & new_n10212_;
  assign new_n10214_ = ~new_n10211_ & new_n10213_;
  assign new_n10215_ = ~new_n4069_ & new_n10122_;
  assign new_n10216_ = new_n10214_ & ~new_n10215_;
  assign new_n10217_ = new_n3820_ & new_n10128_;
  assign new_n10218_ = new_n3870_ & new_n10143_;
  assign new_n10219_ = ~new_n10217_ & ~new_n10218_;
  assign new_n10220_ = new_n10216_ & new_n10219_;
  assign new_n10221_ = ~new_n5105_ & new_n10128_;
  assign new_n10222_ = new_n10220_ & ~new_n10221_;
  assign new_n10223_ = new_n3815_ & new_n10134_;
  assign new_n10224_ = new_n4088_ & new_n10122_;
  assign new_n10225_ = ~new_n10223_ & ~new_n10224_;
  assign new_n10226_ = new_n10206_ & new_n10222_;
  assign new_n10227_ = new_n10225_ & new_n10226_;
  assign new_n10228_ = ~new_n3841_ & new_n10227_;
  assign li0083 = ~new_n10185_ | ~new_n10228_;
  assign new_n10230_ = lo0084 & ~new_n5134_;
  assign new_n10231_ = ~lo0024 & lo0084;
  assign new_n10232_ = new_n4050_ & new_n10231_;
  assign new_n10233_ = lo0084 & new_n5562_;
  assign new_n10234_ = lo0084 & ~lo0314;
  assign new_n10235_ = lo0084 & new_n5155_;
  assign new_n10236_ = new_n3777_ & new_n10235_;
  assign new_n10237_ = lo0084 & ~new_n4632_;
  assign new_n10238_ = new_n5565_ & new_n10237_;
  assign new_n10239_ = ~new_n10236_ & ~new_n10238_;
  assign new_n10240_ = ~new_n5460_ & new_n10234_;
  assign new_n10241_ = new_n10239_ & ~new_n10240_;
  assign new_n10242_ = lo0084 & ~lo0841;
  assign new_n10243_ = new_n3763_ & new_n10242_;
  assign new_n10244_ = new_n3780_ & new_n10231_;
  assign new_n10245_ = ~new_n10243_ & ~new_n10244_;
  assign new_n10246_ = new_n3794_ & new_n10234_;
  assign new_n10247_ = new_n10245_ & ~new_n10246_;
  assign new_n10248_ = ~new_n10232_ & ~new_n10233_;
  assign new_n10249_ = new_n10241_ & new_n10248_;
  assign new_n10250_ = new_n10247_ & new_n10249_;
  assign new_n10251_ = new_n4041_ & new_n10231_;
  assign new_n10252_ = new_n10250_ & ~new_n10251_;
  assign new_n10253_ = new_n3786_ & new_n10231_;
  assign new_n10254_ = lo0084 & new_n5140_;
  assign new_n10255_ = ~new_n10253_ & ~new_n10254_;
  assign new_n10256_ = ~lo1044 & new_n10234_;
  assign new_n10257_ = new_n4007_ & new_n10256_;
  assign new_n10258_ = new_n3969_ & new_n10242_;
  assign new_n10259_ = ~new_n10257_ & ~new_n10258_;
  assign new_n10260_ = new_n3948_ & new_n10231_;
  assign new_n10261_ = new_n10252_ & new_n10255_;
  assign new_n10262_ = new_n10259_ & new_n10261_;
  assign new_n10263_ = ~new_n10260_ & new_n10262_;
  assign new_n10264_ = new_n5133_ & new_n10230_;
  assign new_n10265_ = new_n10263_ & ~new_n10264_;
  assign new_n10266_ = lo0084 & new_n4001_;
  assign new_n10267_ = new_n5230_ & new_n10266_;
  assign new_n10268_ = lo0084 & ~new_n5216_;
  assign new_n10269_ = new_n4133_ & new_n10231_;
  assign new_n10270_ = ~new_n10268_ & ~new_n10269_;
  assign new_n10271_ = lo0084 & li0583;
  assign new_n10272_ = new_n3974_ & new_n10271_;
  assign new_n10273_ = ~new_n4135_ & new_n10272_;
  assign new_n10274_ = lo0084 & new_n5225_;
  assign new_n10275_ = ~new_n10273_ & ~new_n10274_;
  assign new_n10276_ = ~new_n5060_ & new_n10234_;
  assign new_n10277_ = new_n3940_ & new_n10231_;
  assign new_n10278_ = ~new_n10276_ & ~new_n10277_;
  assign new_n10279_ = lo0084 & ~lo0993;
  assign new_n10280_ = new_n3927_ & new_n10279_;
  assign new_n10281_ = new_n3953_ & new_n10231_;
  assign new_n10282_ = ~new_n10280_ & ~new_n10281_;
  assign new_n10283_ = new_n10270_ & new_n10275_;
  assign new_n10284_ = new_n10278_ & new_n10283_;
  assign new_n10285_ = new_n10282_ & new_n10284_;
  assign new_n10286_ = ~new_n5201_ & new_n10242_;
  assign new_n10287_ = lo0084 & new_n5194_;
  assign new_n10288_ = ~new_n10231_ & ~new_n10287_;
  assign new_n10289_ = new_n3936_ & ~new_n10288_;
  assign new_n10290_ = new_n3625_ & new_n10231_;
  assign new_n10291_ = ~new_n10289_ & ~new_n10290_;
  assign new_n10292_ = lo0084 & new_n5818_;
  assign new_n10293_ = ~new_n5184_ & new_n10292_;
  assign new_n10294_ = lo0084 & new_n3706_;
  assign new_n10295_ = ~new_n10286_ & new_n10291_;
  assign new_n10296_ = ~new_n10293_ & new_n10295_;
  assign new_n10297_ = ~new_n10294_ & new_n10296_;
  assign new_n10298_ = new_n10285_ & new_n10297_;
  assign new_n10299_ = new_n10265_ & ~new_n10267_;
  assign new_n10300_ = new_n10298_ & new_n10299_;
  assign new_n10301_ = new_n3804_ & new_n10231_;
  assign new_n10302_ = new_n3834_ & new_n10271_;
  assign new_n10303_ = new_n3678_ & new_n10302_;
  assign new_n10304_ = lo0084 & new_n5112_;
  assign new_n10305_ = new_n3810_ & new_n10242_;
  assign new_n10306_ = ~new_n10301_ & ~new_n10303_;
  assign new_n10307_ = ~new_n10304_ & new_n10306_;
  assign new_n10308_ = ~new_n10305_ & new_n10307_;
  assign new_n10309_ = ~new_n5105_ & new_n10242_;
  assign new_n10310_ = new_n10308_ & ~new_n10309_;
  assign new_n10311_ = new_n3815_ & new_n10234_;
  assign new_n10312_ = new_n4088_ & new_n10231_;
  assign new_n10313_ = ~new_n10311_ & ~new_n10312_;
  assign new_n10314_ = new_n3820_ & new_n10242_;
  assign new_n10315_ = new_n3870_ & new_n10256_;
  assign new_n10316_ = ~new_n10314_ & ~new_n10315_;
  assign new_n10317_ = ~new_n4069_ & new_n10231_;
  assign new_n10318_ = new_n10310_ & new_n10313_;
  assign new_n10319_ = new_n10316_ & new_n10318_;
  assign new_n10320_ = ~new_n10317_ & new_n10319_;
  assign new_n10321_ = new_n4020_ & new_n10231_;
  assign new_n10322_ = ~new_n5096_ & new_n10242_;
  assign new_n10323_ = ~new_n10321_ & ~new_n10322_;
  assign new_n10324_ = lo0314 & new_n6074_;
  assign new_n10325_ = ~new_n10234_ & ~new_n10324_;
  assign new_n10326_ = new_n3746_ & ~new_n10325_;
  assign new_n10327_ = lo0084 & new_n5071_;
  assign new_n10328_ = lo0084 & lo0786;
  assign new_n10329_ = ~new_n5076_ & new_n10271_;
  assign new_n10330_ = lo0084 & new_n5545_;
  assign new_n10331_ = ~new_n10329_ & ~new_n10330_;
  assign new_n10332_ = new_n4475_ & ~new_n10331_;
  assign new_n10333_ = new_n5082_ & new_n10328_;
  assign new_n10334_ = ~new_n10332_ & ~new_n10333_;
  assign new_n10335_ = ~new_n10327_ & new_n10334_;
  assign new_n10336_ = new_n4653_ & ~new_n10335_;
  assign new_n10337_ = ~new_n4096_ & new_n10231_;
  assign new_n10338_ = lo0084 & ~new_n10231_;
  assign new_n10339_ = ~new_n10337_ & ~new_n10338_;
  assign new_n10340_ = new_n4424_ & new_n10336_;
  assign new_n10341_ = new_n5090_ & ~new_n10339_;
  assign new_n10342_ = ~new_n10340_ & ~new_n10341_;
  assign new_n10343_ = new_n10320_ & new_n10323_;
  assign new_n10344_ = ~new_n10326_ & new_n10343_;
  assign new_n10345_ = new_n10342_ & new_n10344_;
  assign li0084 = ~new_n10300_ | ~new_n10345_;
  assign new_n10347_ = ~lo0024 & lo0085;
  assign new_n10348_ = lo0085 & ~lo0841;
  assign new_n10349_ = lo0085 & ~new_n4632_;
  assign new_n10350_ = new_n5565_ & new_n10349_;
  assign new_n10351_ = new_n3763_ & new_n10348_;
  assign new_n10352_ = ~new_n10350_ & ~new_n10351_;
  assign new_n10353_ = lo0085 & ~lo0314;
  assign new_n10354_ = lo0085 & new_n5155_;
  assign new_n10355_ = new_n3903_ & new_n10353_;
  assign new_n10356_ = new_n3777_ & new_n10354_;
  assign new_n10357_ = ~new_n10355_ & ~new_n10356_;
  assign new_n10358_ = lo0085 & new_n5562_;
  assign new_n10359_ = new_n4050_ & new_n10347_;
  assign new_n10360_ = ~new_n10358_ & ~new_n10359_;
  assign new_n10361_ = new_n3780_ & new_n10347_;
  assign new_n10362_ = ~new_n3898_ & new_n10357_;
  assign new_n10363_ = new_n10360_ & new_n10362_;
  assign new_n10364_ = ~new_n10361_ & new_n10363_;
  assign new_n10365_ = ~new_n4575_ & new_n10353_;
  assign new_n10366_ = new_n10364_ & ~new_n10365_;
  assign new_n10367_ = new_n10352_ & new_n10366_;
  assign new_n10368_ = new_n4041_ & new_n10347_;
  assign new_n10369_ = new_n10367_ & ~new_n10368_;
  assign new_n10370_ = new_n3786_ & new_n10347_;
  assign new_n10371_ = lo0085 & new_n5140_;
  assign new_n10372_ = new_n10369_ & ~new_n10370_;
  assign new_n10373_ = ~new_n10371_ & new_n10372_;
  assign new_n10374_ = ~lo1044 & new_n10353_;
  assign new_n10375_ = new_n4007_ & new_n10374_;
  assign new_n10376_ = new_n3969_ & new_n10348_;
  assign new_n10377_ = ~new_n10375_ & ~new_n10376_;
  assign new_n10378_ = new_n3948_ & new_n10347_;
  assign new_n10379_ = lo0085 & li0583;
  assign new_n10380_ = new_n3974_ & new_n10379_;
  assign new_n10381_ = ~new_n4135_ & new_n10380_;
  assign new_n10382_ = lo0085 & new_n5225_;
  assign new_n10383_ = ~new_n10381_ & ~new_n10382_;
  assign new_n10384_ = lo0085 & ~new_n5216_;
  assign new_n10385_ = new_n4133_ & new_n10347_;
  assign new_n10386_ = ~new_n10384_ & ~new_n10385_;
  assign new_n10387_ = new_n10377_ & ~new_n10378_;
  assign new_n10388_ = new_n10383_ & new_n10387_;
  assign new_n10389_ = new_n10386_ & new_n10388_;
  assign new_n10390_ = new_n10373_ & new_n10389_;
  assign new_n10391_ = ~new_n5060_ & new_n10353_;
  assign new_n10392_ = new_n3940_ & new_n10347_;
  assign new_n10393_ = ~new_n10391_ & ~new_n10392_;
  assign new_n10394_ = lo0085 & ~lo0993;
  assign new_n10395_ = new_n3927_ & new_n10394_;
  assign new_n10396_ = new_n3953_ & new_n10347_;
  assign new_n10397_ = ~new_n10395_ & ~new_n10396_;
  assign new_n10398_ = new_n10393_ & new_n10397_;
  assign new_n10399_ = lo0085 & ~new_n5134_;
  assign new_n10400_ = ~new_n5201_ & new_n10348_;
  assign new_n10401_ = lo0085 & new_n5194_;
  assign new_n10402_ = ~new_n10347_ & ~new_n10401_;
  assign new_n10403_ = new_n3936_ & ~new_n10402_;
  assign new_n10404_ = new_n3625_ & new_n10347_;
  assign new_n10405_ = ~new_n10403_ & ~new_n10404_;
  assign new_n10406_ = lo0085 & new_n7163_;
  assign new_n10407_ = lo0085 & new_n3706_;
  assign new_n10408_ = ~new_n10400_ & new_n10405_;
  assign new_n10409_ = ~new_n10406_ & new_n10408_;
  assign new_n10410_ = ~new_n10407_ & new_n10409_;
  assign new_n10411_ = new_n5133_ & new_n10399_;
  assign new_n10412_ = new_n10410_ & ~new_n10411_;
  assign new_n10413_ = lo0085 & new_n5505_;
  assign new_n10414_ = new_n10390_ & new_n10398_;
  assign new_n10415_ = new_n10412_ & new_n10414_;
  assign new_n10416_ = ~new_n10413_ & new_n10415_;
  assign new_n10417_ = new_n3804_ & new_n10347_;
  assign new_n10418_ = new_n3834_ & new_n10379_;
  assign new_n10419_ = new_n3678_ & new_n10418_;
  assign new_n10420_ = lo0085 & new_n5112_;
  assign new_n10421_ = new_n3810_ & new_n10348_;
  assign new_n10422_ = ~new_n10417_ & ~new_n10419_;
  assign new_n10423_ = ~new_n10420_ & new_n10422_;
  assign new_n10424_ = ~new_n10421_ & new_n10423_;
  assign new_n10425_ = ~new_n5105_ & new_n10348_;
  assign new_n10426_ = new_n10424_ & ~new_n10425_;
  assign new_n10427_ = new_n3815_ & new_n10353_;
  assign new_n10428_ = new_n4088_ & new_n10347_;
  assign new_n10429_ = ~new_n10427_ & ~new_n10428_;
  assign new_n10430_ = new_n3820_ & new_n10348_;
  assign new_n10431_ = new_n3870_ & new_n10374_;
  assign new_n10432_ = ~new_n10430_ & ~new_n10431_;
  assign new_n10433_ = ~new_n4069_ & new_n10347_;
  assign new_n10434_ = new_n10426_ & new_n10429_;
  assign new_n10435_ = new_n10432_ & new_n10434_;
  assign new_n10436_ = ~new_n10433_ & new_n10435_;
  assign new_n10437_ = new_n4020_ & new_n10347_;
  assign new_n10438_ = ~new_n5096_ & new_n10348_;
  assign new_n10439_ = ~new_n10437_ & ~new_n10438_;
  assign new_n10440_ = ~new_n4096_ & new_n10347_;
  assign new_n10441_ = lo0085 & ~new_n10347_;
  assign new_n10442_ = ~new_n10440_ & ~new_n10441_;
  assign new_n10443_ = new_n5090_ & ~new_n10442_;
  assign new_n10444_ = new_n3746_ & new_n10353_;
  assign new_n10445_ = ~new_n10443_ & ~new_n10444_;
  assign new_n10446_ = lo0085 & new_n5071_;
  assign new_n10447_ = lo0085 & new_n4219_;
  assign new_n10448_ = ~new_n5074_ & new_n10447_;
  assign new_n10449_ = ~new_n5076_ & new_n10379_;
  assign new_n10450_ = ~new_n10448_ & ~new_n10449_;
  assign new_n10451_ = new_n4475_ & ~new_n10450_;
  assign new_n10452_ = lo0085 & new_n5083_;
  assign new_n10453_ = ~new_n10446_ & ~new_n10451_;
  assign new_n10454_ = ~new_n10452_ & new_n10453_;
  assign new_n10455_ = new_n5070_ & ~new_n10454_;
  assign new_n10456_ = new_n10436_ & new_n10439_;
  assign new_n10457_ = new_n10445_ & new_n10456_;
  assign new_n10458_ = ~new_n10455_ & new_n10457_;
  assign li0085 = ~new_n10416_ | ~new_n10458_;
  assign new_n10460_ = lo0086 & ~lo0841;
  assign new_n10461_ = lo0086 & ~lo0314;
  assign new_n10462_ = ~lo1044 & new_n10461_;
  assign new_n10463_ = new_n4007_ & new_n10462_;
  assign new_n10464_ = new_n3969_ & new_n10460_;
  assign new_n10465_ = ~new_n10463_ & ~new_n10464_;
  assign new_n10466_ = ~lo0024 & lo0086;
  assign new_n10467_ = new_n3786_ & new_n10466_;
  assign new_n10468_ = lo0086 & new_n5140_;
  assign new_n10469_ = new_n3948_ & new_n10466_;
  assign new_n10470_ = new_n10465_ & ~new_n10467_;
  assign new_n10471_ = ~new_n10468_ & new_n10470_;
  assign new_n10472_ = ~new_n10469_ & new_n10471_;
  assign new_n10473_ = ~new_n5060_ & new_n10461_;
  assign new_n10474_ = new_n3940_ & new_n10466_;
  assign new_n10475_ = ~new_n10473_ & ~new_n10474_;
  assign new_n10476_ = lo0086 & ~new_n5216_;
  assign new_n10477_ = new_n4133_ & new_n10466_;
  assign new_n10478_ = ~new_n10476_ & ~new_n10477_;
  assign new_n10479_ = lo0086 & li0583;
  assign new_n10480_ = new_n3974_ & new_n10479_;
  assign new_n10481_ = ~new_n4135_ & new_n10480_;
  assign new_n10482_ = lo0086 & new_n5225_;
  assign new_n10483_ = ~new_n10481_ & ~new_n10482_;
  assign new_n10484_ = lo0086 & ~lo0993;
  assign new_n10485_ = new_n3927_ & new_n10484_;
  assign new_n10486_ = new_n3953_ & new_n10466_;
  assign new_n10487_ = ~new_n10485_ & ~new_n10486_;
  assign new_n10488_ = new_n10475_ & new_n10478_;
  assign new_n10489_ = new_n10483_ & new_n10488_;
  assign new_n10490_ = new_n10487_ & new_n10489_;
  assign new_n10491_ = new_n10472_ & new_n10490_;
  assign new_n10492_ = ~new_n5201_ & new_n10460_;
  assign new_n10493_ = lo0086 & new_n5194_;
  assign new_n10494_ = ~new_n10466_ & ~new_n10493_;
  assign new_n10495_ = new_n3936_ & ~new_n10494_;
  assign new_n10496_ = new_n3625_ & new_n10466_;
  assign new_n10497_ = ~new_n10495_ & ~new_n10496_;
  assign new_n10498_ = lo0086 & new_n5818_;
  assign new_n10499_ = ~new_n5184_ & new_n10498_;
  assign new_n10500_ = lo0086 & new_n3706_;
  assign new_n10501_ = ~new_n10492_ & new_n10497_;
  assign new_n10502_ = ~new_n10499_ & new_n10501_;
  assign new_n10503_ = ~new_n10500_ & new_n10502_;
  assign new_n10504_ = new_n10491_ & new_n10503_;
  assign new_n10505_ = lo0086 & new_n4001_;
  assign new_n10506_ = new_n5230_ & new_n10505_;
  assign new_n10507_ = new_n4050_ & new_n10466_;
  assign new_n10508_ = lo0086 & new_n5562_;
  assign new_n10509_ = lo0086 & new_n5155_;
  assign new_n10510_ = new_n3777_ & new_n10509_;
  assign new_n10511_ = lo0086 & ~new_n4632_;
  assign new_n10512_ = new_n5565_ & new_n10511_;
  assign new_n10513_ = ~new_n10510_ & ~new_n10512_;
  assign new_n10514_ = ~new_n5460_ & new_n10461_;
  assign new_n10515_ = new_n10513_ & ~new_n10514_;
  assign new_n10516_ = new_n3763_ & new_n10460_;
  assign new_n10517_ = new_n3780_ & new_n10466_;
  assign new_n10518_ = ~new_n10516_ & ~new_n10517_;
  assign new_n10519_ = new_n3794_ & new_n10461_;
  assign new_n10520_ = new_n10518_ & ~new_n10519_;
  assign new_n10521_ = ~new_n10507_ & ~new_n10508_;
  assign new_n10522_ = new_n10515_ & new_n10521_;
  assign new_n10523_ = new_n10520_ & new_n10522_;
  assign new_n10524_ = new_n4041_ & new_n10466_;
  assign new_n10525_ = new_n10523_ & ~new_n10524_;
  assign new_n10526_ = lo0086 & ~new_n5134_;
  assign new_n10527_ = new_n5133_ & new_n10526_;
  assign new_n10528_ = new_n10504_ & ~new_n10506_;
  assign new_n10529_ = new_n10525_ & new_n10528_;
  assign new_n10530_ = ~new_n10527_ & new_n10529_;
  assign new_n10531_ = new_n3804_ & new_n10466_;
  assign new_n10532_ = new_n3834_ & new_n10479_;
  assign new_n10533_ = new_n3678_ & new_n10532_;
  assign new_n10534_ = lo0086 & new_n5112_;
  assign new_n10535_ = new_n3810_ & new_n10460_;
  assign new_n10536_ = ~new_n10531_ & ~new_n10533_;
  assign new_n10537_ = ~new_n10534_ & new_n10536_;
  assign new_n10538_ = ~new_n10535_ & new_n10537_;
  assign new_n10539_ = ~new_n5105_ & new_n10460_;
  assign new_n10540_ = new_n10538_ & ~new_n10539_;
  assign new_n10541_ = new_n3815_ & new_n10461_;
  assign new_n10542_ = new_n4088_ & new_n10466_;
  assign new_n10543_ = ~new_n10541_ & ~new_n10542_;
  assign new_n10544_ = new_n3820_ & new_n10460_;
  assign new_n10545_ = new_n3870_ & new_n10462_;
  assign new_n10546_ = ~new_n10544_ & ~new_n10545_;
  assign new_n10547_ = ~new_n4069_ & new_n10466_;
  assign new_n10548_ = new_n10540_ & new_n10543_;
  assign new_n10549_ = new_n10546_ & new_n10548_;
  assign new_n10550_ = ~new_n10547_ & new_n10549_;
  assign new_n10551_ = new_n4020_ & new_n10466_;
  assign new_n10552_ = ~new_n5096_ & new_n10460_;
  assign new_n10553_ = ~new_n10551_ & ~new_n10552_;
  assign new_n10554_ = ~new_n4096_ & new_n10466_;
  assign new_n10555_ = lo0086 & ~new_n10466_;
  assign new_n10556_ = ~new_n10554_ & ~new_n10555_;
  assign new_n10557_ = new_n5090_ & ~new_n10556_;
  assign new_n10558_ = new_n3746_ & new_n10461_;
  assign new_n10559_ = ~new_n10557_ & ~new_n10558_;
  assign new_n10560_ = lo0086 & new_n5071_;
  assign new_n10561_ = lo0086 & lo0786;
  assign new_n10562_ = lo0086 & new_n5545_;
  assign new_n10563_ = new_n4135_ & new_n4228_;
  assign new_n10564_ = ~new_n5076_ & new_n10479_;
  assign new_n10565_ = ~new_n10563_ & ~new_n10564_;
  assign new_n10566_ = ~new_n10562_ & new_n10565_;
  assign new_n10567_ = new_n4475_ & ~new_n10566_;
  assign new_n10568_ = new_n5082_ & new_n10561_;
  assign new_n10569_ = ~new_n10567_ & ~new_n10568_;
  assign new_n10570_ = ~new_n10560_ & new_n10569_;
  assign new_n10571_ = new_n5070_ & ~new_n10570_;
  assign new_n10572_ = new_n10550_ & new_n10553_;
  assign new_n10573_ = new_n10559_ & new_n10572_;
  assign new_n10574_ = ~new_n10571_ & new_n10573_;
  assign li0086 = ~new_n10530_ | ~new_n10574_;
  assign new_n10576_ = ~lo0024 & lo0087;
  assign new_n10577_ = lo0087 & ~lo0314;
  assign new_n10578_ = lo0087 & new_n5155_;
  assign new_n10579_ = new_n3777_ & new_n10578_;
  assign new_n10580_ = lo0087 & ~new_n4632_;
  assign new_n10581_ = new_n5565_ & new_n10580_;
  assign new_n10582_ = ~new_n10579_ & ~new_n10581_;
  assign new_n10583_ = ~new_n5460_ & new_n10577_;
  assign new_n10584_ = new_n10582_ & ~new_n10583_;
  assign new_n10585_ = lo0087 & new_n5562_;
  assign new_n10586_ = new_n4050_ & new_n10576_;
  assign new_n10587_ = lo0087 & ~lo0841;
  assign new_n10588_ = new_n3763_ & new_n10587_;
  assign new_n10589_ = new_n3780_ & new_n10576_;
  assign new_n10590_ = ~new_n10588_ & ~new_n10589_;
  assign new_n10591_ = new_n3794_ & new_n10577_;
  assign new_n10592_ = new_n10590_ & ~new_n10591_;
  assign new_n10593_ = new_n10584_ & ~new_n10585_;
  assign new_n10594_ = ~new_n10586_ & new_n10593_;
  assign new_n10595_ = new_n10592_ & new_n10594_;
  assign new_n10596_ = new_n4041_ & new_n10576_;
  assign new_n10597_ = new_n10595_ & ~new_n10596_;
  assign new_n10598_ = lo0087 & new_n3678_;
  assign new_n10599_ = new_n3786_ & new_n10576_;
  assign new_n10600_ = new_n5139_ & new_n10598_;
  assign new_n10601_ = ~new_n10599_ & ~new_n10600_;
  assign new_n10602_ = ~lo1044 & new_n10577_;
  assign new_n10603_ = new_n4007_ & new_n10602_;
  assign new_n10604_ = new_n3969_ & new_n10587_;
  assign new_n10605_ = ~new_n10603_ & ~new_n10604_;
  assign new_n10606_ = lo0087 & ~new_n5216_;
  assign new_n10607_ = new_n4133_ & new_n10576_;
  assign new_n10608_ = ~new_n10606_ & ~new_n10607_;
  assign new_n10609_ = lo0087 & li0583;
  assign new_n10610_ = new_n3974_ & new_n10609_;
  assign new_n10611_ = ~new_n4135_ & new_n10610_;
  assign new_n10612_ = lo0087 & new_n5225_;
  assign new_n10613_ = new_n10608_ & ~new_n10611_;
  assign new_n10614_ = ~new_n10612_ & new_n10613_;
  assign new_n10615_ = new_n3948_ & new_n10576_;
  assign new_n10616_ = new_n10614_ & ~new_n10615_;
  assign new_n10617_ = new_n10597_ & new_n10601_;
  assign new_n10618_ = new_n10605_ & new_n10617_;
  assign new_n10619_ = new_n10616_ & new_n10618_;
  assign new_n10620_ = lo0087 & new_n5505_;
  assign new_n10621_ = lo0087 & new_n5135_;
  assign new_n10622_ = lo0087 & new_n5194_;
  assign new_n10623_ = ~new_n10576_ & ~new_n10622_;
  assign new_n10624_ = new_n3936_ & ~new_n10623_;
  assign new_n10625_ = new_n3625_ & new_n10576_;
  assign new_n10626_ = ~new_n10624_ & ~new_n10625_;
  assign new_n10627_ = lo0087 & new_n3706_;
  assign new_n10628_ = lo0087 & new_n5708_;
  assign new_n10629_ = new_n10626_ & ~new_n10627_;
  assign new_n10630_ = ~new_n10628_ & new_n10629_;
  assign new_n10631_ = ~new_n5201_ & new_n10587_;
  assign new_n10632_ = new_n10630_ & ~new_n10631_;
  assign new_n10633_ = ~new_n10620_ & ~new_n10621_;
  assign new_n10634_ = new_n10632_ & new_n10633_;
  assign new_n10635_ = new_n10619_ & new_n10634_;
  assign new_n10636_ = ~new_n5105_ & new_n10587_;
  assign new_n10637_ = ~new_n5060_ & new_n10577_;
  assign new_n10638_ = new_n3940_ & new_n10576_;
  assign new_n10639_ = ~new_n10637_ & ~new_n10638_;
  assign new_n10640_ = lo0087 & ~lo0993;
  assign new_n10641_ = new_n3927_ & new_n10640_;
  assign new_n10642_ = new_n3953_ & new_n10576_;
  assign new_n10643_ = ~new_n10641_ & ~new_n10642_;
  assign new_n10644_ = new_n10639_ & new_n10643_;
  assign new_n10645_ = new_n4020_ & new_n10576_;
  assign new_n10646_ = ~new_n5096_ & new_n10587_;
  assign new_n10647_ = ~new_n10645_ & ~new_n10646_;
  assign new_n10648_ = lo0087 & new_n5071_;
  assign new_n10649_ = lo0087 & new_n4219_;
  assign new_n10650_ = ~new_n5074_ & new_n10649_;
  assign new_n10651_ = ~new_n5076_ & new_n10609_;
  assign new_n10652_ = ~new_n10650_ & ~new_n10651_;
  assign new_n10653_ = new_n4475_ & ~new_n10652_;
  assign new_n10654_ = lo0087 & new_n5083_;
  assign new_n10655_ = ~new_n10648_ & ~new_n10653_;
  assign new_n10656_ = ~new_n10654_ & new_n10655_;
  assign new_n10657_ = new_n5070_ & ~new_n10656_;
  assign new_n10658_ = ~new_n4096_ & new_n10576_;
  assign new_n10659_ = lo0087 & ~new_n10576_;
  assign new_n10660_ = ~new_n10658_ & ~new_n10659_;
  assign new_n10661_ = new_n5090_ & ~new_n10660_;
  assign new_n10662_ = new_n3746_ & new_n10577_;
  assign new_n10663_ = ~new_n10661_ & ~new_n10662_;
  assign new_n10664_ = new_n10647_ & ~new_n10657_;
  assign new_n10665_ = new_n10663_ & new_n10664_;
  assign new_n10666_ = ~lo0087 & ~lo0314;
  assign new_n10667_ = new_n3815_ & ~new_n10666_;
  assign new_n10668_ = new_n3804_ & new_n10576_;
  assign new_n10669_ = new_n3834_ & new_n10609_;
  assign new_n10670_ = new_n3678_ & new_n10669_;
  assign new_n10671_ = lo0087 & new_n5112_;
  assign new_n10672_ = new_n3810_ & new_n10587_;
  assign new_n10673_ = ~new_n10668_ & ~new_n10670_;
  assign new_n10674_ = ~new_n10671_ & new_n10673_;
  assign new_n10675_ = ~new_n10672_ & new_n10674_;
  assign new_n10676_ = new_n4088_ & new_n10576_;
  assign new_n10677_ = new_n10675_ & ~new_n10676_;
  assign new_n10678_ = new_n3820_ & new_n10587_;
  assign new_n10679_ = new_n3870_ & new_n10602_;
  assign new_n10680_ = ~new_n10678_ & ~new_n10679_;
  assign new_n10681_ = ~new_n4069_ & new_n10576_;
  assign new_n10682_ = ~new_n10667_ & new_n10677_;
  assign new_n10683_ = new_n10680_ & new_n10682_;
  assign new_n10684_ = ~new_n10681_ & new_n10683_;
  assign new_n10685_ = new_n10665_ & new_n10684_;
  assign new_n10686_ = new_n10635_ & ~new_n10636_;
  assign new_n10687_ = new_n10644_ & new_n10686_;
  assign li0087 = ~new_n10685_ | ~new_n10687_;
  assign new_n10689_ = lo0088 & ~lo0841;
  assign new_n10690_ = ~lo0024 & lo0088;
  assign new_n10691_ = new_n3804_ & new_n10690_;
  assign new_n10692_ = lo0088 & li0583;
  assign new_n10693_ = new_n3834_ & new_n10692_;
  assign new_n10694_ = new_n3678_ & new_n10693_;
  assign new_n10695_ = lo0088 & new_n5112_;
  assign new_n10696_ = new_n3810_ & new_n10689_;
  assign new_n10697_ = ~new_n10691_ & ~new_n10694_;
  assign new_n10698_ = ~new_n10695_ & new_n10697_;
  assign new_n10699_ = ~new_n10696_ & new_n10698_;
  assign new_n10700_ = ~new_n5105_ & new_n10689_;
  assign new_n10701_ = new_n10699_ & ~new_n10700_;
  assign new_n10702_ = lo0088 & ~lo0314;
  assign new_n10703_ = new_n3815_ & new_n10702_;
  assign new_n10704_ = new_n4088_ & new_n10690_;
  assign new_n10705_ = ~new_n10703_ & ~new_n10704_;
  assign new_n10706_ = ~lo1044 & new_n10702_;
  assign new_n10707_ = new_n3820_ & new_n10689_;
  assign new_n10708_ = new_n3870_ & new_n10706_;
  assign new_n10709_ = ~new_n10707_ & ~new_n10708_;
  assign new_n10710_ = ~new_n4069_ & new_n10690_;
  assign new_n10711_ = new_n10701_ & new_n10705_;
  assign new_n10712_ = new_n10709_ & new_n10711_;
  assign new_n10713_ = ~new_n10710_ & new_n10712_;
  assign new_n10714_ = lo0088 & new_n3678_;
  assign new_n10715_ = ~new_n5137_ & ~new_n10714_;
  assign new_n10716_ = new_n3891_ & ~new_n10715_;
  assign new_n10717_ = lo0088 & new_n5562_;
  assign new_n10718_ = lo0088 & new_n5155_;
  assign new_n10719_ = new_n3777_ & new_n10718_;
  assign new_n10720_ = lo0088 & ~new_n4632_;
  assign new_n10721_ = new_n5565_ & new_n10720_;
  assign new_n10722_ = ~new_n10719_ & ~new_n10721_;
  assign new_n10723_ = ~new_n5460_ & new_n10702_;
  assign new_n10724_ = new_n10722_ & ~new_n10723_;
  assign new_n10725_ = new_n3763_ & new_n10689_;
  assign new_n10726_ = new_n3780_ & new_n10690_;
  assign new_n10727_ = ~new_n10725_ & ~new_n10726_;
  assign new_n10728_ = new_n3794_ & new_n10702_;
  assign new_n10729_ = new_n10727_ & ~new_n10728_;
  assign new_n10730_ = ~new_n10716_ & ~new_n10717_;
  assign new_n10731_ = new_n10724_ & new_n10730_;
  assign new_n10732_ = new_n10729_ & new_n10731_;
  assign new_n10733_ = ~new_n6390_ & new_n10690_;
  assign new_n10734_ = new_n10732_ & ~new_n10733_;
  assign new_n10735_ = lo0088 & ~new_n5216_;
  assign new_n10736_ = new_n4133_ & new_n10690_;
  assign new_n10737_ = ~new_n10735_ & ~new_n10736_;
  assign new_n10738_ = new_n3974_ & new_n10692_;
  assign new_n10739_ = ~new_n4135_ & new_n10738_;
  assign new_n10740_ = lo0088 & new_n5225_;
  assign new_n10741_ = new_n10737_ & ~new_n10739_;
  assign new_n10742_ = ~new_n10740_ & new_n10741_;
  assign new_n10743_ = new_n3948_ & new_n10690_;
  assign new_n10744_ = new_n10742_ & ~new_n10743_;
  assign new_n10745_ = new_n4007_ & new_n10706_;
  assign new_n10746_ = new_n3969_ & new_n10689_;
  assign new_n10747_ = ~new_n10745_ & ~new_n10746_;
  assign new_n10748_ = new_n10734_ & new_n10744_;
  assign new_n10749_ = new_n10747_ & new_n10748_;
  assign new_n10750_ = lo0088 & new_n5071_;
  assign new_n10751_ = lo0088 & new_n4219_;
  assign new_n10752_ = ~new_n5074_ & new_n10751_;
  assign new_n10753_ = ~new_n5076_ & new_n10692_;
  assign new_n10754_ = ~new_n10752_ & ~new_n10753_;
  assign new_n10755_ = new_n4475_ & ~new_n10754_;
  assign new_n10756_ = lo0088 & new_n5083_;
  assign new_n10757_ = ~new_n10750_ & ~new_n10755_;
  assign new_n10758_ = ~new_n10756_ & new_n10757_;
  assign new_n10759_ = new_n5070_ & ~new_n10758_;
  assign new_n10760_ = ~new_n4096_ & new_n10690_;
  assign new_n10761_ = lo0088 & ~new_n10690_;
  assign new_n10762_ = ~new_n10760_ & ~new_n10761_;
  assign new_n10763_ = new_n5090_ & ~new_n10762_;
  assign new_n10764_ = new_n3746_ & new_n10702_;
  assign new_n10765_ = ~new_n10763_ & ~new_n10764_;
  assign new_n10766_ = new_n4020_ & new_n10690_;
  assign new_n10767_ = ~new_n5096_ & new_n10689_;
  assign new_n10768_ = ~new_n10766_ & ~new_n10767_;
  assign new_n10769_ = ~new_n10759_ & new_n10765_;
  assign new_n10770_ = new_n10768_ & new_n10769_;
  assign new_n10771_ = new_n10749_ & new_n10770_;
  assign new_n10772_ = lo0088 & new_n5505_;
  assign new_n10773_ = lo0088 & ~new_n5134_;
  assign new_n10774_ = new_n5133_ & new_n10773_;
  assign new_n10775_ = ~new_n5060_ & new_n10702_;
  assign new_n10776_ = new_n3940_ & new_n10690_;
  assign new_n10777_ = ~new_n10775_ & ~new_n10776_;
  assign new_n10778_ = lo0088 & ~lo0993;
  assign new_n10779_ = new_n3927_ & new_n10778_;
  assign new_n10780_ = new_n3953_ & new_n10690_;
  assign new_n10781_ = ~new_n10779_ & ~new_n10780_;
  assign new_n10782_ = ~new_n10772_ & ~new_n10774_;
  assign new_n10783_ = new_n10777_ & new_n10782_;
  assign new_n10784_ = new_n10781_ & new_n10783_;
  assign new_n10785_ = ~new_n5201_ & new_n10689_;
  assign new_n10786_ = lo0088 & new_n5194_;
  assign new_n10787_ = ~new_n10690_ & ~new_n10786_;
  assign new_n10788_ = new_n3936_ & ~new_n10787_;
  assign new_n10789_ = new_n3625_ & new_n10690_;
  assign new_n10790_ = ~new_n10788_ & ~new_n10789_;
  assign new_n10791_ = lo0088 & new_n5608_;
  assign new_n10792_ = ~new_n5184_ & new_n10791_;
  assign new_n10793_ = lo0088 & new_n3706_;
  assign new_n10794_ = ~new_n10785_ & new_n10790_;
  assign new_n10795_ = ~new_n10792_ & new_n10794_;
  assign new_n10796_ = ~new_n10793_ & new_n10795_;
  assign new_n10797_ = new_n10784_ & new_n10796_;
  assign new_n10798_ = new_n10713_ & new_n10771_;
  assign li0088 = ~new_n10797_ | ~new_n10798_;
  assign new_n10800_ = lo0089 & ~new_n5134_;
  assign new_n10801_ = new_n5133_ & new_n10800_;
  assign new_n10802_ = lo0089 & li0583;
  assign new_n10803_ = new_n3974_ & new_n10802_;
  assign new_n10804_ = ~new_n4135_ & new_n10803_;
  assign new_n10805_ = lo0089 & new_n5225_;
  assign new_n10806_ = ~new_n10804_ & ~new_n10805_;
  assign new_n10807_ = lo0089 & ~lo0841;
  assign new_n10808_ = lo0089 & ~lo0314;
  assign new_n10809_ = ~lo1044 & new_n10808_;
  assign new_n10810_ = new_n4007_ & new_n10809_;
  assign new_n10811_ = new_n3969_ & new_n10807_;
  assign new_n10812_ = ~new_n10810_ & ~new_n10811_;
  assign new_n10813_ = ~lo0024 & lo0089;
  assign new_n10814_ = new_n3948_ & new_n10813_;
  assign new_n10815_ = ~new_n10801_ & new_n10806_;
  assign new_n10816_ = new_n10812_ & new_n10815_;
  assign new_n10817_ = ~new_n10814_ & new_n10816_;
  assign new_n10818_ = ~new_n5201_ & new_n10807_;
  assign new_n10819_ = lo0089 & new_n5194_;
  assign new_n10820_ = ~new_n10813_ & ~new_n10819_;
  assign new_n10821_ = new_n3936_ & ~new_n10820_;
  assign new_n10822_ = new_n3625_ & new_n10813_;
  assign new_n10823_ = ~new_n10821_ & ~new_n10822_;
  assign new_n10824_ = lo0089 & new_n5608_;
  assign new_n10825_ = ~new_n5184_ & new_n10824_;
  assign new_n10826_ = lo0089 & new_n3706_;
  assign new_n10827_ = ~new_n10818_ & new_n10823_;
  assign new_n10828_ = ~new_n10825_ & new_n10827_;
  assign new_n10829_ = ~new_n10826_ & new_n10828_;
  assign new_n10830_ = new_n10817_ & new_n10829_;
  assign new_n10831_ = new_n4050_ & new_n10813_;
  assign new_n10832_ = lo0089 & new_n5562_;
  assign new_n10833_ = lo0089 & new_n5155_;
  assign new_n10834_ = new_n3777_ & new_n10833_;
  assign new_n10835_ = lo0089 & ~new_n4632_;
  assign new_n10836_ = new_n5565_ & new_n10835_;
  assign new_n10837_ = ~new_n10834_ & ~new_n10836_;
  assign new_n10838_ = ~new_n5460_ & new_n10808_;
  assign new_n10839_ = new_n10837_ & ~new_n10838_;
  assign new_n10840_ = new_n3763_ & new_n10807_;
  assign new_n10841_ = new_n3780_ & new_n10813_;
  assign new_n10842_ = ~new_n10840_ & ~new_n10841_;
  assign new_n10843_ = new_n3794_ & new_n10808_;
  assign new_n10844_ = new_n10842_ & ~new_n10843_;
  assign new_n10845_ = ~new_n10831_ & ~new_n10832_;
  assign new_n10846_ = new_n10839_ & new_n10845_;
  assign new_n10847_ = new_n10844_ & new_n10846_;
  assign new_n10848_ = new_n4041_ & new_n10813_;
  assign new_n10849_ = new_n10847_ & ~new_n10848_;
  assign new_n10850_ = lo0089 & new_n4001_;
  assign new_n10851_ = new_n5230_ & new_n10850_;
  assign new_n10852_ = ~new_n5060_ & new_n10808_;
  assign new_n10853_ = new_n3940_ & new_n10813_;
  assign new_n10854_ = ~new_n10852_ & ~new_n10853_;
  assign new_n10855_ = lo0089 & ~lo0993;
  assign new_n10856_ = new_n3927_ & new_n10855_;
  assign new_n10857_ = new_n3953_ & new_n10813_;
  assign new_n10858_ = ~new_n10856_ & ~new_n10857_;
  assign new_n10859_ = new_n10854_ & new_n10858_;
  assign new_n10860_ = lo0089 & ~new_n5216_;
  assign new_n10861_ = new_n4133_ & new_n10813_;
  assign new_n10862_ = ~new_n10860_ & ~new_n10861_;
  assign new_n10863_ = new_n3786_ & new_n10813_;
  assign new_n10864_ = lo0089 & new_n5140_;
  assign new_n10865_ = new_n10862_ & ~new_n10863_;
  assign new_n10866_ = ~new_n10864_ & new_n10865_;
  assign new_n10867_ = new_n10859_ & new_n10866_;
  assign new_n10868_ = new_n10830_ & new_n10849_;
  assign new_n10869_ = ~new_n10851_ & new_n10868_;
  assign new_n10870_ = new_n10867_ & new_n10869_;
  assign new_n10871_ = lo0089 & new_n5112_;
  assign new_n10872_ = new_n3810_ & new_n10807_;
  assign new_n10873_ = new_n3834_ & new_n10802_;
  assign new_n10874_ = new_n3678_ & new_n10873_;
  assign new_n10875_ = ~lo0024 & ~lo0089;
  assign new_n10876_ = new_n3804_ & ~new_n10875_;
  assign new_n10877_ = ~new_n10871_ & ~new_n10872_;
  assign new_n10878_ = ~new_n10874_ & new_n10877_;
  assign new_n10879_ = ~new_n10876_ & new_n10878_;
  assign new_n10880_ = ~new_n5105_ & new_n10807_;
  assign new_n10881_ = new_n10879_ & ~new_n10880_;
  assign new_n10882_ = new_n3815_ & new_n10808_;
  assign new_n10883_ = new_n4088_ & new_n10813_;
  assign new_n10884_ = ~new_n10882_ & ~new_n10883_;
  assign new_n10885_ = new_n3820_ & new_n10807_;
  assign new_n10886_ = new_n3870_ & new_n10809_;
  assign new_n10887_ = ~new_n10885_ & ~new_n10886_;
  assign new_n10888_ = ~new_n4069_ & new_n10813_;
  assign new_n10889_ = new_n10881_ & new_n10884_;
  assign new_n10890_ = new_n10887_ & new_n10889_;
  assign new_n10891_ = ~new_n10888_ & new_n10890_;
  assign new_n10892_ = new_n4020_ & new_n10813_;
  assign new_n10893_ = ~new_n5096_ & new_n10807_;
  assign new_n10894_ = ~new_n10892_ & ~new_n10893_;
  assign new_n10895_ = ~new_n4096_ & new_n10813_;
  assign new_n10896_ = lo0089 & ~new_n10813_;
  assign new_n10897_ = ~new_n10895_ & ~new_n10896_;
  assign new_n10898_ = new_n5090_ & ~new_n10897_;
  assign new_n10899_ = new_n3746_ & new_n10808_;
  assign new_n10900_ = ~new_n10898_ & ~new_n10899_;
  assign new_n10901_ = lo0089 & new_n5071_;
  assign new_n10902_ = lo0089 & new_n4219_;
  assign new_n10903_ = ~new_n5074_ & new_n10902_;
  assign new_n10904_ = ~new_n5076_ & new_n10802_;
  assign new_n10905_ = ~new_n10903_ & ~new_n10904_;
  assign new_n10906_ = new_n4475_ & ~new_n10905_;
  assign new_n10907_ = lo0089 & new_n5083_;
  assign new_n10908_ = ~new_n10901_ & ~new_n10906_;
  assign new_n10909_ = ~new_n10907_ & new_n10908_;
  assign new_n10910_ = new_n5070_ & ~new_n10909_;
  assign new_n10911_ = new_n10891_ & new_n10894_;
  assign new_n10912_ = new_n10900_ & new_n10911_;
  assign new_n10913_ = ~new_n10910_ & new_n10912_;
  assign li0089 = ~new_n10870_ | ~new_n10913_;
  assign new_n10915_ = lo0090 & ~lo0314;
  assign new_n10916_ = ~lo0024 & lo0090;
  assign new_n10917_ = ~new_n5060_ & new_n10915_;
  assign new_n10918_ = new_n3940_ & new_n10916_;
  assign new_n10919_ = ~new_n10917_ & ~new_n10918_;
  assign new_n10920_ = lo0090 & ~lo0993;
  assign new_n10921_ = new_n3927_ & new_n10920_;
  assign new_n10922_ = new_n3953_ & new_n10916_;
  assign new_n10923_ = ~new_n10921_ & ~new_n10922_;
  assign new_n10924_ = new_n10919_ & new_n10923_;
  assign new_n10925_ = new_n4050_ & new_n10916_;
  assign new_n10926_ = new_n3794_ & new_n10915_;
  assign new_n10927_ = lo0090 & new_n3773_;
  assign new_n10928_ = lo1076 & new_n10927_;
  assign new_n10929_ = ~new_n5460_ & new_n10915_;
  assign new_n10930_ = ~new_n10925_ & ~new_n10926_;
  assign new_n10931_ = ~new_n10928_ & new_n10930_;
  assign new_n10932_ = ~new_n10929_ & new_n10931_;
  assign new_n10933_ = lo0090 & ~lo0841;
  assign new_n10934_ = new_n3763_ & new_n10933_;
  assign new_n10935_ = new_n3780_ & new_n10916_;
  assign new_n10936_ = ~new_n10934_ & ~new_n10935_;
  assign new_n10937_ = new_n10932_ & new_n10936_;
  assign new_n10938_ = lo0090 & ~new_n4632_;
  assign new_n10939_ = lo0090 & new_n5155_;
  assign new_n10940_ = new_n3777_ & new_n10939_;
  assign new_n10941_ = new_n5565_ & new_n10938_;
  assign new_n10942_ = ~new_n10940_ & ~new_n10941_;
  assign new_n10943_ = new_n10937_ & new_n10942_;
  assign new_n10944_ = new_n4041_ & new_n10916_;
  assign new_n10945_ = new_n10943_ & ~new_n10944_;
  assign new_n10946_ = new_n3786_ & new_n10916_;
  assign new_n10947_ = lo0090 & new_n5140_;
  assign new_n10948_ = new_n10945_ & ~new_n10946_;
  assign new_n10949_ = ~new_n10947_ & new_n10948_;
  assign new_n10950_ = new_n3969_ & new_n10933_;
  assign new_n10951_ = new_n4007_ & new_n10915_;
  assign new_n10952_ = ~lo1044 & new_n10951_;
  assign new_n10953_ = ~new_n10950_ & ~new_n10952_;
  assign new_n10954_ = new_n3948_ & new_n10916_;
  assign new_n10955_ = new_n10953_ & ~new_n10954_;
  assign new_n10956_ = lo0090 & ~new_n5216_;
  assign new_n10957_ = new_n4133_ & new_n10916_;
  assign new_n10958_ = ~new_n10956_ & ~new_n10957_;
  assign new_n10959_ = lo0090 & new_n5225_;
  assign new_n10960_ = lo0090 & li0583;
  assign new_n10961_ = new_n3974_ & new_n10960_;
  assign new_n10962_ = ~new_n4135_ & new_n10961_;
  assign new_n10963_ = new_n10955_ & new_n10958_;
  assign new_n10964_ = ~new_n10959_ & new_n10963_;
  assign new_n10965_ = ~new_n10962_ & new_n10964_;
  assign new_n10966_ = new_n10949_ & new_n10965_;
  assign new_n10967_ = lo0090 & ~new_n5134_;
  assign new_n10968_ = ~new_n5201_ & new_n10933_;
  assign new_n10969_ = lo0090 & new_n5194_;
  assign new_n10970_ = ~new_n10916_ & ~new_n10969_;
  assign new_n10971_ = new_n3936_ & ~new_n10970_;
  assign new_n10972_ = new_n3625_ & new_n10916_;
  assign new_n10973_ = ~new_n10971_ & ~new_n10972_;
  assign new_n10974_ = lo0090 & new_n5608_;
  assign new_n10975_ = ~new_n5184_ & new_n10974_;
  assign new_n10976_ = lo0090 & new_n3706_;
  assign new_n10977_ = ~new_n10968_ & new_n10973_;
  assign new_n10978_ = ~new_n10975_ & new_n10977_;
  assign new_n10979_ = ~new_n10976_ & new_n10978_;
  assign new_n10980_ = new_n5133_ & new_n10967_;
  assign new_n10981_ = new_n10979_ & ~new_n10980_;
  assign new_n10982_ = lo0090 & new_n5505_;
  assign new_n10983_ = new_n10924_ & new_n10966_;
  assign new_n10984_ = new_n10981_ & new_n10983_;
  assign new_n10985_ = ~new_n10982_ & new_n10984_;
  assign new_n10986_ = ~new_n5096_ & new_n10933_;
  assign new_n10987_ = new_n4020_ & new_n10916_;
  assign new_n10988_ = ~new_n10986_ & ~new_n10987_;
  assign new_n10989_ = lo0090 & new_n5071_;
  assign new_n10990_ = lo0090 & lo0786;
  assign new_n10991_ = ~new_n5076_ & new_n10960_;
  assign new_n10992_ = lo0090 & new_n5545_;
  assign new_n10993_ = ~new_n10991_ & ~new_n10992_;
  assign new_n10994_ = new_n4475_ & ~new_n10993_;
  assign new_n10995_ = new_n5082_ & new_n10990_;
  assign new_n10996_ = ~new_n10994_ & ~new_n10995_;
  assign new_n10997_ = ~new_n10989_ & new_n10996_;
  assign new_n10998_ = new_n5070_ & ~new_n10997_;
  assign new_n10999_ = new_n3746_ & new_n10915_;
  assign new_n11000_ = ~new_n4096_ & new_n10916_;
  assign new_n11001_ = lo0090 & ~new_n10916_;
  assign new_n11002_ = ~new_n11000_ & ~new_n11001_;
  assign new_n11003_ = new_n5090_ & ~new_n11002_;
  assign new_n11004_ = ~new_n10999_ & ~new_n11003_;
  assign new_n11005_ = ~new_n10998_ & new_n11004_;
  assign new_n11006_ = new_n10988_ & new_n11005_;
  assign new_n11007_ = lo0090 & new_n5112_;
  assign new_n11008_ = new_n3810_ & new_n10933_;
  assign new_n11009_ = new_n3834_ & new_n10960_;
  assign new_n11010_ = new_n3678_ & new_n11009_;
  assign new_n11011_ = ~lo1044 & ~new_n10915_;
  assign new_n11012_ = new_n3870_ & ~new_n11011_;
  assign new_n11013_ = ~new_n11007_ & ~new_n11008_;
  assign new_n11014_ = ~new_n11010_ & new_n11013_;
  assign new_n11015_ = ~new_n11012_ & new_n11014_;
  assign new_n11016_ = ~new_n5105_ & new_n10933_;
  assign new_n11017_ = new_n11015_ & ~new_n11016_;
  assign new_n11018_ = new_n3815_ & new_n10915_;
  assign new_n11019_ = new_n4088_ & new_n10916_;
  assign new_n11020_ = ~new_n11018_ & ~new_n11019_;
  assign new_n11021_ = new_n3820_ & new_n10933_;
  assign new_n11022_ = new_n3618_ & new_n10916_;
  assign new_n11023_ = ~new_n11021_ & ~new_n11022_;
  assign new_n11024_ = ~new_n5394_ & new_n10916_;
  assign new_n11025_ = new_n11023_ & ~new_n11024_;
  assign new_n11026_ = new_n11006_ & new_n11017_;
  assign new_n11027_ = new_n11020_ & new_n11026_;
  assign new_n11028_ = new_n11025_ & new_n11027_;
  assign li0090 = ~new_n10985_ | ~new_n11028_;
  assign new_n11030_ = lo0091 & ~lo0314;
  assign new_n11031_ = ~lo0024 & lo0091;
  assign new_n11032_ = ~new_n5060_ & new_n11030_;
  assign new_n11033_ = new_n3940_ & new_n11031_;
  assign new_n11034_ = ~new_n11032_ & ~new_n11033_;
  assign new_n11035_ = lo0091 & ~lo0993;
  assign new_n11036_ = new_n3927_ & new_n11035_;
  assign new_n11037_ = new_n3953_ & new_n11031_;
  assign new_n11038_ = ~new_n11036_ & ~new_n11037_;
  assign new_n11039_ = new_n11034_ & new_n11038_;
  assign new_n11040_ = new_n4050_ & new_n11031_;
  assign new_n11041_ = lo0091 & new_n5562_;
  assign new_n11042_ = lo0091 & new_n5155_;
  assign new_n11043_ = new_n3777_ & new_n11042_;
  assign new_n11044_ = lo0091 & ~new_n4632_;
  assign new_n11045_ = new_n5565_ & new_n11044_;
  assign new_n11046_ = ~new_n11043_ & ~new_n11045_;
  assign new_n11047_ = ~new_n5460_ & new_n11030_;
  assign new_n11048_ = new_n11046_ & ~new_n11047_;
  assign new_n11049_ = lo0091 & ~lo0841;
  assign new_n11050_ = new_n3763_ & new_n11049_;
  assign new_n11051_ = new_n3780_ & new_n11031_;
  assign new_n11052_ = ~new_n11050_ & ~new_n11051_;
  assign new_n11053_ = new_n3794_ & new_n11030_;
  assign new_n11054_ = new_n11052_ & ~new_n11053_;
  assign new_n11055_ = ~new_n11040_ & ~new_n11041_;
  assign new_n11056_ = new_n11048_ & new_n11055_;
  assign new_n11057_ = new_n11054_ & new_n11056_;
  assign new_n11058_ = new_n4041_ & new_n11031_;
  assign new_n11059_ = new_n11057_ & ~new_n11058_;
  assign new_n11060_ = new_n3786_ & new_n11031_;
  assign new_n11061_ = lo0091 & new_n5140_;
  assign new_n11062_ = new_n11059_ & ~new_n11060_;
  assign new_n11063_ = ~new_n11061_ & new_n11062_;
  assign new_n11064_ = ~lo1044 & new_n11030_;
  assign new_n11065_ = new_n4007_ & new_n11064_;
  assign new_n11066_ = new_n3969_ & new_n11049_;
  assign new_n11067_ = ~new_n11065_ & ~new_n11066_;
  assign new_n11068_ = new_n3948_ & new_n11031_;
  assign new_n11069_ = lo0091 & li0583;
  assign new_n11070_ = new_n3974_ & new_n11069_;
  assign new_n11071_ = ~new_n4135_ & new_n11070_;
  assign new_n11072_ = lo0091 & new_n5225_;
  assign new_n11073_ = ~new_n11071_ & ~new_n11072_;
  assign new_n11074_ = lo0091 & ~new_n5216_;
  assign new_n11075_ = new_n4133_ & new_n11031_;
  assign new_n11076_ = ~new_n11074_ & ~new_n11075_;
  assign new_n11077_ = new_n11067_ & ~new_n11068_;
  assign new_n11078_ = new_n11073_ & new_n11077_;
  assign new_n11079_ = new_n11076_ & new_n11078_;
  assign new_n11080_ = new_n11063_ & new_n11079_;
  assign new_n11081_ = lo0091 & ~new_n5134_;
  assign new_n11082_ = ~new_n5201_ & new_n11049_;
  assign new_n11083_ = lo0091 & new_n5194_;
  assign new_n11084_ = ~new_n11031_ & ~new_n11083_;
  assign new_n11085_ = new_n3936_ & ~new_n11084_;
  assign new_n11086_ = new_n3625_ & new_n11031_;
  assign new_n11087_ = ~new_n11085_ & ~new_n11086_;
  assign new_n11088_ = lo0091 & new_n5818_;
  assign new_n11089_ = ~new_n5184_ & new_n11088_;
  assign new_n11090_ = lo0091 & new_n3706_;
  assign new_n11091_ = ~new_n11082_ & new_n11087_;
  assign new_n11092_ = ~new_n11089_ & new_n11091_;
  assign new_n11093_ = ~new_n11090_ & new_n11092_;
  assign new_n11094_ = new_n5133_ & new_n11081_;
  assign new_n11095_ = new_n11093_ & ~new_n11094_;
  assign new_n11096_ = lo0091 & new_n5505_;
  assign new_n11097_ = new_n11039_ & new_n11080_;
  assign new_n11098_ = new_n11095_ & new_n11097_;
  assign new_n11099_ = ~new_n11096_ & new_n11098_;
  assign new_n11100_ = new_n3804_ & new_n11031_;
  assign new_n11101_ = new_n3834_ & new_n11069_;
  assign new_n11102_ = new_n3678_ & new_n11101_;
  assign new_n11103_ = lo0091 & new_n5112_;
  assign new_n11104_ = new_n3810_ & new_n11049_;
  assign new_n11105_ = ~new_n11100_ & ~new_n11102_;
  assign new_n11106_ = ~new_n11103_ & new_n11105_;
  assign new_n11107_ = ~new_n11104_ & new_n11106_;
  assign new_n11108_ = ~new_n5105_ & new_n11049_;
  assign new_n11109_ = new_n11107_ & ~new_n11108_;
  assign new_n11110_ = new_n3815_ & new_n11030_;
  assign new_n11111_ = new_n4088_ & new_n11031_;
  assign new_n11112_ = ~new_n11110_ & ~new_n11111_;
  assign new_n11113_ = new_n3820_ & new_n11049_;
  assign new_n11114_ = new_n3870_ & new_n11064_;
  assign new_n11115_ = ~new_n11113_ & ~new_n11114_;
  assign new_n11116_ = ~new_n4069_ & new_n11031_;
  assign new_n11117_ = new_n11109_ & new_n11112_;
  assign new_n11118_ = new_n11115_ & new_n11117_;
  assign new_n11119_ = ~new_n11116_ & new_n11118_;
  assign new_n11120_ = new_n3746_ & new_n11030_;
  assign new_n11121_ = new_n4020_ & new_n11031_;
  assign new_n11122_ = ~new_n11120_ & ~new_n11121_;
  assign new_n11123_ = ~new_n5096_ & new_n11049_;
  assign new_n11124_ = new_n11122_ & ~new_n11123_;
  assign new_n11125_ = new_n3753_ & new_n4135_;
  assign new_n11126_ = lo0091 & new_n5071_;
  assign new_n11127_ = lo0091 & lo0786;
  assign new_n11128_ = lo0091 & new_n5545_;
  assign new_n11129_ = ~new_n5076_ & new_n11069_;
  assign new_n11130_ = ~new_n4655_ & ~new_n11129_;
  assign new_n11131_ = ~new_n11128_ & new_n11130_;
  assign new_n11132_ = new_n4475_ & ~new_n11131_;
  assign new_n11133_ = new_n5082_ & new_n11127_;
  assign new_n11134_ = ~new_n11132_ & ~new_n11133_;
  assign new_n11135_ = ~new_n11126_ & new_n11134_;
  assign new_n11136_ = new_n4653_ & ~new_n11135_;
  assign new_n11137_ = ~new_n4096_ & new_n11031_;
  assign new_n11138_ = lo0091 & ~new_n11031_;
  assign new_n11139_ = ~new_n11137_ & ~new_n11138_;
  assign new_n11140_ = new_n4424_ & new_n11136_;
  assign new_n11141_ = new_n5090_ & ~new_n11139_;
  assign new_n11142_ = ~new_n11140_ & ~new_n11141_;
  assign new_n11143_ = new_n11119_ & new_n11124_;
  assign new_n11144_ = ~new_n11125_ & new_n11143_;
  assign new_n11145_ = new_n11142_ & new_n11144_;
  assign li0091 = ~new_n11099_ | ~new_n11145_;
  assign new_n11147_ = lo0092 & ~new_n5134_;
  assign new_n11148_ = new_n5133_ & new_n11147_;
  assign new_n11149_ = lo0092 & li0583;
  assign new_n11150_ = new_n3974_ & new_n11149_;
  assign new_n11151_ = ~new_n4135_ & new_n11150_;
  assign new_n11152_ = lo0092 & new_n5225_;
  assign new_n11153_ = ~new_n11151_ & ~new_n11152_;
  assign new_n11154_ = lo0092 & ~lo0841;
  assign new_n11155_ = lo0092 & ~lo0314;
  assign new_n11156_ = ~lo1044 & new_n11155_;
  assign new_n11157_ = new_n4007_ & new_n11156_;
  assign new_n11158_ = new_n3969_ & new_n11154_;
  assign new_n11159_ = ~new_n11157_ & ~new_n11158_;
  assign new_n11160_ = ~lo0024 & lo0092;
  assign new_n11161_ = new_n3948_ & new_n11160_;
  assign new_n11162_ = ~new_n11148_ & new_n11153_;
  assign new_n11163_ = new_n11159_ & new_n11162_;
  assign new_n11164_ = ~new_n11161_ & new_n11163_;
  assign new_n11165_ = ~new_n5201_ & new_n11154_;
  assign new_n11166_ = lo0092 & new_n5194_;
  assign new_n11167_ = ~new_n11160_ & ~new_n11166_;
  assign new_n11168_ = new_n3936_ & ~new_n11167_;
  assign new_n11169_ = new_n3625_ & new_n11160_;
  assign new_n11170_ = ~new_n11168_ & ~new_n11169_;
  assign new_n11171_ = lo0092 & new_n5818_;
  assign new_n11172_ = ~new_n5184_ & new_n11171_;
  assign new_n11173_ = lo0092 & new_n3706_;
  assign new_n11174_ = ~new_n11165_ & new_n11170_;
  assign new_n11175_ = ~new_n11172_ & new_n11174_;
  assign new_n11176_ = ~new_n11173_ & new_n11175_;
  assign new_n11177_ = new_n11164_ & new_n11176_;
  assign new_n11178_ = new_n4050_ & new_n11160_;
  assign new_n11179_ = lo0092 & new_n5562_;
  assign new_n11180_ = lo0092 & new_n5155_;
  assign new_n11181_ = new_n3777_ & new_n11180_;
  assign new_n11182_ = lo0092 & ~new_n4632_;
  assign new_n11183_ = new_n5565_ & new_n11182_;
  assign new_n11184_ = ~new_n11181_ & ~new_n11183_;
  assign new_n11185_ = ~new_n5460_ & new_n11155_;
  assign new_n11186_ = new_n11184_ & ~new_n11185_;
  assign new_n11187_ = new_n3763_ & new_n11154_;
  assign new_n11188_ = new_n3780_ & new_n11160_;
  assign new_n11189_ = ~new_n11187_ & ~new_n11188_;
  assign new_n11190_ = new_n3794_ & new_n11155_;
  assign new_n11191_ = new_n11189_ & ~new_n11190_;
  assign new_n11192_ = ~new_n11178_ & ~new_n11179_;
  assign new_n11193_ = new_n11186_ & new_n11192_;
  assign new_n11194_ = new_n11191_ & new_n11193_;
  assign new_n11195_ = new_n4041_ & new_n11160_;
  assign new_n11196_ = new_n11194_ & ~new_n11195_;
  assign new_n11197_ = lo0092 & new_n4001_;
  assign new_n11198_ = new_n5230_ & new_n11197_;
  assign new_n11199_ = ~new_n5060_ & new_n11155_;
  assign new_n11200_ = new_n3940_ & new_n11160_;
  assign new_n11201_ = ~new_n11199_ & ~new_n11200_;
  assign new_n11202_ = lo0092 & ~lo0993;
  assign new_n11203_ = new_n3927_ & new_n11202_;
  assign new_n11204_ = new_n3953_ & new_n11160_;
  assign new_n11205_ = ~new_n11203_ & ~new_n11204_;
  assign new_n11206_ = new_n11201_ & new_n11205_;
  assign new_n11207_ = lo0092 & ~new_n5216_;
  assign new_n11208_ = new_n4133_ & new_n11160_;
  assign new_n11209_ = ~new_n11207_ & ~new_n11208_;
  assign new_n11210_ = new_n3786_ & new_n11160_;
  assign new_n11211_ = lo0092 & new_n5140_;
  assign new_n11212_ = new_n11209_ & ~new_n11210_;
  assign new_n11213_ = ~new_n11211_ & new_n11212_;
  assign new_n11214_ = new_n11206_ & new_n11213_;
  assign new_n11215_ = new_n11177_ & new_n11196_;
  assign new_n11216_ = ~new_n11198_ & new_n11215_;
  assign new_n11217_ = new_n11214_ & new_n11216_;
  assign new_n11218_ = new_n3804_ & new_n11160_;
  assign new_n11219_ = new_n3834_ & new_n11149_;
  assign new_n11220_ = new_n3678_ & new_n11219_;
  assign new_n11221_ = lo0092 & new_n5112_;
  assign new_n11222_ = new_n3810_ & new_n11154_;
  assign new_n11223_ = ~new_n11218_ & ~new_n11220_;
  assign new_n11224_ = ~new_n11221_ & new_n11223_;
  assign new_n11225_ = ~new_n11222_ & new_n11224_;
  assign new_n11226_ = ~new_n5105_ & new_n11154_;
  assign new_n11227_ = new_n11225_ & ~new_n11226_;
  assign new_n11228_ = new_n3815_ & new_n11155_;
  assign new_n11229_ = new_n4088_ & new_n11160_;
  assign new_n11230_ = ~new_n11228_ & ~new_n11229_;
  assign new_n11231_ = new_n3820_ & new_n11154_;
  assign new_n11232_ = new_n3870_ & new_n11156_;
  assign new_n11233_ = ~new_n11231_ & ~new_n11232_;
  assign new_n11234_ = ~new_n4069_ & new_n11160_;
  assign new_n11235_ = new_n11227_ & new_n11230_;
  assign new_n11236_ = new_n11233_ & new_n11235_;
  assign new_n11237_ = ~new_n11234_ & new_n11236_;
  assign new_n11238_ = new_n4020_ & new_n11160_;
  assign new_n11239_ = ~new_n5096_ & new_n11154_;
  assign new_n11240_ = ~new_n11238_ & ~new_n11239_;
  assign new_n11241_ = ~new_n4096_ & new_n11160_;
  assign new_n11242_ = lo0092 & ~new_n11160_;
  assign new_n11243_ = ~new_n11241_ & ~new_n11242_;
  assign new_n11244_ = new_n5090_ & ~new_n11243_;
  assign new_n11245_ = new_n3746_ & new_n11155_;
  assign new_n11246_ = ~new_n11244_ & ~new_n11245_;
  assign new_n11247_ = lo0092 & new_n5071_;
  assign new_n11248_ = lo0092 & lo0786;
  assign new_n11249_ = lo0092 & new_n5545_;
  assign new_n11250_ = new_n4135_ & new_n4428_;
  assign new_n11251_ = ~new_n5076_ & new_n11149_;
  assign new_n11252_ = ~new_n11250_ & ~new_n11251_;
  assign new_n11253_ = ~new_n11249_ & new_n11252_;
  assign new_n11254_ = new_n4475_ & ~new_n11253_;
  assign new_n11255_ = new_n5082_ & new_n11248_;
  assign new_n11256_ = ~new_n11254_ & ~new_n11255_;
  assign new_n11257_ = ~new_n11247_ & new_n11256_;
  assign new_n11258_ = new_n5070_ & ~new_n11257_;
  assign new_n11259_ = new_n11237_ & new_n11240_;
  assign new_n11260_ = new_n11246_ & new_n11259_;
  assign new_n11261_ = ~new_n11258_ & new_n11260_;
  assign li0092 = ~new_n11217_ | ~new_n11261_;
  assign new_n11263_ = lo0093 & ~lo0314;
  assign new_n11264_ = ~lo0024 & lo0093;
  assign new_n11265_ = ~new_n5060_ & new_n11263_;
  assign new_n11266_ = new_n3940_ & new_n11264_;
  assign new_n11267_ = ~new_n11265_ & ~new_n11266_;
  assign new_n11268_ = lo0093 & ~lo0993;
  assign new_n11269_ = new_n3927_ & new_n11268_;
  assign new_n11270_ = new_n3953_ & new_n11264_;
  assign new_n11271_ = ~new_n11269_ & ~new_n11270_;
  assign new_n11272_ = new_n11267_ & new_n11271_;
  assign new_n11273_ = new_n4050_ & new_n11264_;
  assign new_n11274_ = lo0093 & new_n5562_;
  assign new_n11275_ = lo0093 & new_n5155_;
  assign new_n11276_ = new_n3777_ & new_n11275_;
  assign new_n11277_ = lo0093 & ~new_n4632_;
  assign new_n11278_ = new_n5565_ & new_n11277_;
  assign new_n11279_ = ~new_n11276_ & ~new_n11278_;
  assign new_n11280_ = ~new_n5460_ & new_n11263_;
  assign new_n11281_ = new_n11279_ & ~new_n11280_;
  assign new_n11282_ = lo0093 & ~lo0841;
  assign new_n11283_ = new_n3763_ & new_n11282_;
  assign new_n11284_ = new_n3780_ & new_n11264_;
  assign new_n11285_ = ~new_n11283_ & ~new_n11284_;
  assign new_n11286_ = new_n3794_ & new_n11263_;
  assign new_n11287_ = new_n11285_ & ~new_n11286_;
  assign new_n11288_ = ~new_n11273_ & ~new_n11274_;
  assign new_n11289_ = new_n11281_ & new_n11288_;
  assign new_n11290_ = new_n11287_ & new_n11289_;
  assign new_n11291_ = new_n4041_ & new_n11264_;
  assign new_n11292_ = new_n11290_ & ~new_n11291_;
  assign new_n11293_ = new_n3786_ & new_n11264_;
  assign new_n11294_ = lo0093 & new_n5140_;
  assign new_n11295_ = new_n11292_ & ~new_n11293_;
  assign new_n11296_ = ~new_n11294_ & new_n11295_;
  assign new_n11297_ = new_n3969_ & new_n11282_;
  assign new_n11298_ = new_n3948_ & new_n11264_;
  assign new_n11299_ = ~new_n11297_ & ~new_n11298_;
  assign new_n11300_ = new_n4133_ & new_n11264_;
  assign new_n11301_ = ~lo1044 & ~new_n11263_;
  assign new_n11302_ = new_n4007_ & ~new_n11301_;
  assign new_n11303_ = lo0093 & li0583;
  assign new_n11304_ = ~new_n4135_ & new_n11303_;
  assign new_n11305_ = new_n3974_ & new_n11304_;
  assign new_n11306_ = lo0093 & ~new_n4135_;
  assign new_n11307_ = new_n5224_ & new_n11306_;
  assign new_n11308_ = ~new_n11305_ & ~new_n11307_;
  assign new_n11309_ = ~new_n11302_ & new_n11308_;
  assign new_n11310_ = lo0093 & ~new_n5216_;
  assign new_n11311_ = new_n11299_ & ~new_n11300_;
  assign new_n11312_ = new_n11309_ & new_n11311_;
  assign new_n11313_ = ~new_n11310_ & new_n11312_;
  assign new_n11314_ = new_n11296_ & new_n11313_;
  assign new_n11315_ = lo0093 & ~new_n5134_;
  assign new_n11316_ = ~new_n5201_ & new_n11282_;
  assign new_n11317_ = lo0093 & new_n5194_;
  assign new_n11318_ = ~new_n11264_ & ~new_n11317_;
  assign new_n11319_ = new_n3936_ & ~new_n11318_;
  assign new_n11320_ = new_n3625_ & new_n11264_;
  assign new_n11321_ = ~new_n11319_ & ~new_n11320_;
  assign new_n11322_ = lo0093 & new_n5818_;
  assign new_n11323_ = ~new_n5184_ & new_n11322_;
  assign new_n11324_ = lo0093 & new_n3706_;
  assign new_n11325_ = ~new_n11316_ & new_n11321_;
  assign new_n11326_ = ~new_n11323_ & new_n11325_;
  assign new_n11327_ = ~new_n11324_ & new_n11326_;
  assign new_n11328_ = new_n5133_ & new_n11315_;
  assign new_n11329_ = new_n11327_ & ~new_n11328_;
  assign new_n11330_ = lo0093 & new_n5505_;
  assign new_n11331_ = new_n11272_ & new_n11314_;
  assign new_n11332_ = new_n11329_ & new_n11331_;
  assign new_n11333_ = ~new_n11330_ & new_n11332_;
  assign new_n11334_ = ~new_n5096_ & new_n11282_;
  assign new_n11335_ = new_n4020_ & new_n11264_;
  assign new_n11336_ = ~new_n11334_ & ~new_n11335_;
  assign new_n11337_ = lo0093 & new_n5071_;
  assign new_n11338_ = lo0093 & lo0786;
  assign new_n11339_ = ~new_n5076_ & new_n11303_;
  assign new_n11340_ = lo0093 & new_n5545_;
  assign new_n11341_ = ~new_n11339_ & ~new_n11340_;
  assign new_n11342_ = new_n4475_ & ~new_n11341_;
  assign new_n11343_ = new_n5082_ & new_n11338_;
  assign new_n11344_ = ~new_n11342_ & ~new_n11343_;
  assign new_n11345_ = ~new_n11337_ & new_n11344_;
  assign new_n11346_ = new_n5070_ & ~new_n11345_;
  assign new_n11347_ = new_n3746_ & new_n11263_;
  assign new_n11348_ = ~new_n4096_ & new_n11264_;
  assign new_n11349_ = lo0093 & ~new_n11264_;
  assign new_n11350_ = ~new_n11348_ & ~new_n11349_;
  assign new_n11351_ = new_n5090_ & ~new_n11350_;
  assign new_n11352_ = ~new_n11347_ & ~new_n11351_;
  assign new_n11353_ = ~new_n11346_ & new_n11352_;
  assign new_n11354_ = new_n11336_ & new_n11353_;
  assign new_n11355_ = new_n3804_ & new_n11264_;
  assign new_n11356_ = new_n3834_ & new_n11303_;
  assign new_n11357_ = new_n3678_ & new_n11356_;
  assign new_n11358_ = lo0093 & new_n5112_;
  assign new_n11359_ = new_n3810_ & new_n11282_;
  assign new_n11360_ = ~new_n11355_ & ~new_n11357_;
  assign new_n11361_ = ~new_n11358_ & new_n11360_;
  assign new_n11362_ = ~new_n11359_ & new_n11361_;
  assign new_n11363_ = ~new_n5105_ & new_n11282_;
  assign new_n11364_ = new_n11362_ & ~new_n11363_;
  assign new_n11365_ = new_n3815_ & new_n11263_;
  assign new_n11366_ = new_n4088_ & new_n11264_;
  assign new_n11367_ = ~new_n11365_ & ~new_n11366_;
  assign new_n11368_ = new_n3820_ & new_n11282_;
  assign new_n11369_ = new_n3870_ & new_n11263_;
  assign new_n11370_ = ~lo1044 & new_n11369_;
  assign new_n11371_ = ~new_n11368_ & ~new_n11370_;
  assign new_n11372_ = ~new_n4069_ & new_n11264_;
  assign new_n11373_ = new_n11371_ & ~new_n11372_;
  assign new_n11374_ = new_n11354_ & new_n11364_;
  assign new_n11375_ = new_n11367_ & new_n11374_;
  assign new_n11376_ = new_n11373_ & new_n11375_;
  assign li0093 = ~new_n11333_ | ~new_n11376_;
  assign new_n11378_ = ~lo0024 & lo0094;
  assign new_n11379_ = lo0094 & ~lo0841;
  assign new_n11380_ = ~new_n5096_ & new_n11379_;
  assign new_n11381_ = new_n4020_ & new_n11378_;
  assign new_n11382_ = ~new_n11380_ & ~new_n11381_;
  assign new_n11383_ = lo0094 & new_n5071_;
  assign new_n11384_ = lo0094 & lo0786;
  assign new_n11385_ = lo0094 & li0583;
  assign new_n11386_ = ~new_n5076_ & new_n11385_;
  assign new_n11387_ = lo0094 & new_n5545_;
  assign new_n11388_ = ~new_n11386_ & ~new_n11387_;
  assign new_n11389_ = new_n4475_ & ~new_n11388_;
  assign new_n11390_ = new_n5082_ & new_n11384_;
  assign new_n11391_ = ~new_n11389_ & ~new_n11390_;
  assign new_n11392_ = ~new_n11383_ & new_n11391_;
  assign new_n11393_ = new_n5070_ & ~new_n11392_;
  assign new_n11394_ = lo0094 & ~lo0314;
  assign new_n11395_ = new_n3746_ & new_n11394_;
  assign new_n11396_ = ~new_n4096_ & new_n11378_;
  assign new_n11397_ = lo0094 & ~new_n11378_;
  assign new_n11398_ = ~new_n11396_ & ~new_n11397_;
  assign new_n11399_ = new_n5090_ & ~new_n11398_;
  assign new_n11400_ = ~new_n11395_ & ~new_n11399_;
  assign new_n11401_ = ~new_n11393_ & new_n11400_;
  assign new_n11402_ = new_n11382_ & new_n11401_;
  assign new_n11403_ = lo0094 & new_n5112_;
  assign new_n11404_ = new_n3810_ & new_n11379_;
  assign new_n11405_ = new_n3834_ & new_n11385_;
  assign new_n11406_ = new_n3678_ & new_n11405_;
  assign new_n11407_ = ~lo0094 & ~lo0841;
  assign new_n11408_ = new_n3820_ & ~new_n11407_;
  assign new_n11409_ = ~new_n11403_ & ~new_n11404_;
  assign new_n11410_ = ~new_n11406_ & new_n11409_;
  assign new_n11411_ = ~new_n11408_ & new_n11410_;
  assign new_n11412_ = ~new_n5105_ & new_n11379_;
  assign new_n11413_ = new_n11411_ & ~new_n11412_;
  assign new_n11414_ = new_n3815_ & new_n11394_;
  assign new_n11415_ = new_n4088_ & new_n11378_;
  assign new_n11416_ = ~new_n11414_ & ~new_n11415_;
  assign new_n11417_ = ~lo1044 & new_n11394_;
  assign new_n11418_ = new_n3618_ & new_n11378_;
  assign new_n11419_ = new_n3870_ & new_n11417_;
  assign new_n11420_ = ~new_n11418_ & ~new_n11419_;
  assign new_n11421_ = ~new_n5394_ & new_n11378_;
  assign new_n11422_ = new_n11420_ & ~new_n11421_;
  assign new_n11423_ = new_n11402_ & new_n11413_;
  assign new_n11424_ = new_n11416_ & new_n11423_;
  assign new_n11425_ = new_n11422_ & new_n11424_;
  assign new_n11426_ = ~new_n5060_ & new_n11394_;
  assign new_n11427_ = new_n3940_ & new_n11378_;
  assign new_n11428_ = ~new_n11426_ & ~new_n11427_;
  assign new_n11429_ = new_n3953_ & new_n11378_;
  assign new_n11430_ = lo0094 & new_n5671_;
  assign new_n11431_ = new_n11428_ & ~new_n11429_;
  assign new_n11432_ = ~new_n11430_ & new_n11431_;
  assign new_n11433_ = lo0094 & new_n5505_;
  assign new_n11434_ = lo0094 & new_n5135_;
  assign new_n11435_ = ~new_n5201_ & new_n11379_;
  assign new_n11436_ = ~new_n11433_ & ~new_n11434_;
  assign new_n11437_ = ~new_n11435_ & new_n11436_;
  assign new_n11438_ = lo0094 & new_n5194_;
  assign new_n11439_ = ~new_n11378_ & ~new_n11438_;
  assign new_n11440_ = new_n3936_ & ~new_n11439_;
  assign new_n11441_ = new_n3625_ & new_n11378_;
  assign new_n11442_ = ~new_n11440_ & ~new_n11441_;
  assign new_n11443_ = lo0094 & new_n3706_;
  assign new_n11444_ = lo0094 & new_n5818_;
  assign new_n11445_ = ~new_n5184_ & new_n11444_;
  assign new_n11446_ = new_n11442_ & ~new_n11443_;
  assign new_n11447_ = ~new_n11445_ & new_n11446_;
  assign new_n11448_ = new_n11437_ & new_n11447_;
  assign new_n11449_ = new_n3786_ & new_n11378_;
  assign new_n11450_ = new_n4007_ & new_n11417_;
  assign new_n11451_ = lo0094 & new_n5562_;
  assign new_n11452_ = new_n4041_ & new_n11378_;
  assign new_n11453_ = ~new_n11450_ & ~new_n11451_;
  assign new_n11454_ = ~new_n11452_ & new_n11453_;
  assign new_n11455_ = ~new_n11449_ & new_n11454_;
  assign new_n11456_ = new_n4050_ & new_n11378_;
  assign new_n11457_ = new_n3969_ & new_n11379_;
  assign new_n11458_ = lo0094 & new_n3678_;
  assign new_n11459_ = new_n5139_ & new_n11458_;
  assign new_n11460_ = new_n3948_ & new_n11378_;
  assign new_n11461_ = ~new_n11459_ & ~new_n11460_;
  assign new_n11462_ = new_n11455_ & ~new_n11456_;
  assign new_n11463_ = ~new_n11457_ & new_n11462_;
  assign new_n11464_ = new_n11461_ & new_n11463_;
  assign new_n11465_ = lo0094 & ~new_n5216_;
  assign new_n11466_ = new_n4133_ & new_n11378_;
  assign new_n11467_ = ~new_n11465_ & ~new_n11466_;
  assign new_n11468_ = new_n3974_ & new_n11385_;
  assign new_n11469_ = ~new_n4135_ & new_n11468_;
  assign new_n11470_ = lo0094 & new_n5225_;
  assign new_n11471_ = new_n11467_ & ~new_n11469_;
  assign new_n11472_ = ~new_n11470_ & new_n11471_;
  assign new_n11473_ = new_n11464_ & new_n11472_;
  assign new_n11474_ = new_n3763_ & new_n11379_;
  assign new_n11475_ = new_n3780_ & new_n11378_;
  assign new_n11476_ = ~new_n11474_ & ~new_n11475_;
  assign new_n11477_ = new_n3794_ & new_n11394_;
  assign new_n11478_ = new_n11476_ & ~new_n11477_;
  assign new_n11479_ = lo0094 & new_n5155_;
  assign new_n11480_ = new_n3777_ & new_n11479_;
  assign new_n11481_ = lo0094 & ~new_n4632_;
  assign new_n11482_ = new_n5565_ & new_n11481_;
  assign new_n11483_ = ~new_n11480_ & ~new_n11482_;
  assign new_n11484_ = ~new_n5460_ & new_n11394_;
  assign new_n11485_ = new_n11483_ & ~new_n11484_;
  assign new_n11486_ = new_n11473_ & new_n11478_;
  assign new_n11487_ = new_n11485_ & new_n11486_;
  assign new_n11488_ = new_n11425_ & new_n11432_;
  assign new_n11489_ = new_n11448_ & new_n11488_;
  assign li0094 = ~new_n11487_ | ~new_n11489_;
  assign new_n11491_ = lo0095 & ~lo0841;
  assign new_n11492_ = ~lo0024 & lo0095;
  assign new_n11493_ = new_n3804_ & new_n11492_;
  assign new_n11494_ = lo0095 & li0583;
  assign new_n11495_ = new_n3834_ & new_n11494_;
  assign new_n11496_ = new_n3678_ & new_n11495_;
  assign new_n11497_ = lo0095 & new_n5112_;
  assign new_n11498_ = new_n3810_ & new_n11491_;
  assign new_n11499_ = ~new_n11493_ & ~new_n11496_;
  assign new_n11500_ = ~new_n11497_ & new_n11499_;
  assign new_n11501_ = ~new_n11498_ & new_n11500_;
  assign new_n11502_ = ~new_n5105_ & new_n11491_;
  assign new_n11503_ = new_n11501_ & ~new_n11502_;
  assign new_n11504_ = lo0095 & ~lo0314;
  assign new_n11505_ = ~lo1044 & new_n11504_;
  assign new_n11506_ = new_n3820_ & new_n11491_;
  assign new_n11507_ = new_n3870_ & new_n11505_;
  assign new_n11508_ = ~new_n11506_ & ~new_n11507_;
  assign new_n11509_ = ~new_n4069_ & new_n11492_;
  assign new_n11510_ = new_n11508_ & ~new_n11509_;
  assign new_n11511_ = new_n3815_ & new_n11504_;
  assign new_n11512_ = new_n4088_ & new_n11492_;
  assign new_n11513_ = ~new_n11511_ & ~new_n11512_;
  assign new_n11514_ = new_n11510_ & new_n11513_;
  assign new_n11515_ = new_n4020_ & new_n11492_;
  assign new_n11516_ = new_n3735_ & new_n11491_;
  assign new_n11517_ = ~new_n11515_ & ~new_n11516_;
  assign new_n11518_ = ~lo0332 & lo0841;
  assign new_n11519_ = ~new_n11491_ & ~new_n11518_;
  assign new_n11520_ = lo0095 & new_n5071_;
  assign new_n11521_ = lo0095 & lo0786;
  assign new_n11522_ = ~new_n8960_ & ~new_n8961_;
  assign new_n11523_ = new_n5074_ & ~new_n11522_;
  assign new_n11524_ = ~lo0095 & ~new_n5074_;
  assign new_n11525_ = ~new_n11523_ & ~new_n11524_;
  assign new_n11526_ = new_n4219_ & new_n11525_;
  assign new_n11527_ = ~new_n5076_ & new_n11494_;
  assign new_n11528_ = ~new_n11526_ & ~new_n11527_;
  assign new_n11529_ = new_n4475_ & ~new_n11528_;
  assign new_n11530_ = new_n5082_ & new_n11521_;
  assign new_n11531_ = ~new_n11529_ & ~new_n11530_;
  assign new_n11532_ = ~new_n11520_ & new_n11531_;
  assign new_n11533_ = new_n4653_ & ~new_n11532_;
  assign new_n11534_ = ~new_n4096_ & new_n11492_;
  assign new_n11535_ = lo0095 & ~new_n11492_;
  assign new_n11536_ = ~new_n11534_ & ~new_n11535_;
  assign new_n11537_ = new_n4424_ & new_n11533_;
  assign new_n11538_ = new_n5090_ & ~new_n11536_;
  assign new_n11539_ = ~new_n11537_ & ~new_n11538_;
  assign new_n11540_ = new_n3589_ & ~new_n11519_;
  assign new_n11541_ = new_n11539_ & ~new_n11540_;
  assign new_n11542_ = new_n3746_ & new_n11504_;
  assign new_n11543_ = new_n11541_ & ~new_n11542_;
  assign new_n11544_ = new_n11503_ & new_n11514_;
  assign new_n11545_ = new_n11517_ & new_n11544_;
  assign new_n11546_ = new_n11543_ & new_n11545_;
  assign new_n11547_ = lo0095 & ~new_n5134_;
  assign new_n11548_ = ~new_n5060_ & new_n11504_;
  assign new_n11549_ = new_n3940_ & new_n11492_;
  assign new_n11550_ = ~new_n11548_ & ~new_n11549_;
  assign new_n11551_ = new_n4007_ & new_n11505_;
  assign new_n11552_ = new_n3969_ & new_n11491_;
  assign new_n11553_ = ~new_n11551_ & ~new_n11552_;
  assign new_n11554_ = lo0095 & ~lo0993;
  assign new_n11555_ = new_n3927_ & new_n11554_;
  assign new_n11556_ = new_n3953_ & new_n11492_;
  assign new_n11557_ = ~new_n11555_ & ~new_n11556_;
  assign new_n11558_ = new_n3948_ & new_n11492_;
  assign new_n11559_ = new_n11550_ & new_n11553_;
  assign new_n11560_ = new_n11557_ & new_n11559_;
  assign new_n11561_ = ~new_n11558_ & new_n11560_;
  assign new_n11562_ = new_n5133_ & new_n11547_;
  assign new_n11563_ = new_n11561_ & ~new_n11562_;
  assign new_n11564_ = ~new_n5201_ & new_n11491_;
  assign new_n11565_ = lo0095 & new_n5194_;
  assign new_n11566_ = ~new_n11492_ & ~new_n11565_;
  assign new_n11567_ = new_n3936_ & ~new_n11566_;
  assign new_n11568_ = new_n3625_ & new_n11492_;
  assign new_n11569_ = ~new_n11567_ & ~new_n11568_;
  assign new_n11570_ = lo0095 & new_n5818_;
  assign new_n11571_ = ~new_n5184_ & new_n11570_;
  assign new_n11572_ = lo0095 & new_n3706_;
  assign new_n11573_ = ~new_n11564_ & new_n11569_;
  assign new_n11574_ = ~new_n11571_ & new_n11573_;
  assign new_n11575_ = ~new_n11572_ & new_n11574_;
  assign new_n11576_ = new_n11563_ & new_n11575_;
  assign new_n11577_ = lo0095 & new_n4001_;
  assign new_n11578_ = new_n5230_ & new_n11577_;
  assign new_n11579_ = new_n4050_ & new_n11492_;
  assign new_n11580_ = lo0095 & new_n5562_;
  assign new_n11581_ = lo0095 & new_n5155_;
  assign new_n11582_ = new_n3777_ & new_n11581_;
  assign new_n11583_ = lo0095 & ~new_n4632_;
  assign new_n11584_ = new_n5565_ & new_n11583_;
  assign new_n11585_ = ~new_n11582_ & ~new_n11584_;
  assign new_n11586_ = ~new_n5460_ & new_n11504_;
  assign new_n11587_ = new_n11585_ & ~new_n11586_;
  assign new_n11588_ = new_n3763_ & new_n11491_;
  assign new_n11589_ = new_n3780_ & new_n11492_;
  assign new_n11590_ = ~new_n11588_ & ~new_n11589_;
  assign new_n11591_ = new_n3794_ & new_n11504_;
  assign new_n11592_ = new_n11590_ & ~new_n11591_;
  assign new_n11593_ = ~new_n11579_ & ~new_n11580_;
  assign new_n11594_ = new_n11587_ & new_n11593_;
  assign new_n11595_ = new_n11592_ & new_n11594_;
  assign new_n11596_ = new_n4041_ & new_n11492_;
  assign new_n11597_ = new_n11595_ & ~new_n11596_;
  assign new_n11598_ = new_n3974_ & new_n11494_;
  assign new_n11599_ = ~new_n4135_ & new_n11598_;
  assign new_n11600_ = lo0095 & new_n5225_;
  assign new_n11601_ = ~new_n11599_ & ~new_n11600_;
  assign new_n11602_ = lo0095 & ~new_n5216_;
  assign new_n11603_ = new_n4133_ & new_n11492_;
  assign new_n11604_ = ~new_n11602_ & ~new_n11603_;
  assign new_n11605_ = new_n3786_ & new_n11492_;
  assign new_n11606_ = lo0095 & new_n5140_;
  assign new_n11607_ = new_n11601_ & new_n11604_;
  assign new_n11608_ = ~new_n11605_ & new_n11607_;
  assign new_n11609_ = ~new_n11606_ & new_n11608_;
  assign new_n11610_ = new_n11576_ & ~new_n11578_;
  assign new_n11611_ = new_n11597_ & new_n11610_;
  assign new_n11612_ = new_n11609_ & new_n11611_;
  assign li0095 = ~new_n11546_ | ~new_n11612_;
  assign new_n11614_ = lo0096 & ~lo0314;
  assign new_n11615_ = ~lo0024 & lo0096;
  assign new_n11616_ = ~new_n5060_ & new_n11614_;
  assign new_n11617_ = new_n3940_ & new_n11615_;
  assign new_n11618_ = ~new_n11616_ & ~new_n11617_;
  assign new_n11619_ = lo0096 & ~lo0993;
  assign new_n11620_ = new_n3927_ & new_n11619_;
  assign new_n11621_ = new_n3953_ & new_n11615_;
  assign new_n11622_ = ~new_n11620_ & ~new_n11621_;
  assign new_n11623_ = new_n11618_ & new_n11622_;
  assign new_n11624_ = new_n4050_ & new_n11615_;
  assign new_n11625_ = lo0096 & new_n5562_;
  assign new_n11626_ = lo0096 & new_n5155_;
  assign new_n11627_ = new_n3777_ & new_n11626_;
  assign new_n11628_ = lo0096 & ~new_n4632_;
  assign new_n11629_ = new_n5565_ & new_n11628_;
  assign new_n11630_ = ~new_n11627_ & ~new_n11629_;
  assign new_n11631_ = ~new_n5460_ & new_n11614_;
  assign new_n11632_ = new_n11630_ & ~new_n11631_;
  assign new_n11633_ = lo0096 & ~lo0841;
  assign new_n11634_ = new_n3763_ & new_n11633_;
  assign new_n11635_ = new_n3780_ & new_n11615_;
  assign new_n11636_ = ~new_n11634_ & ~new_n11635_;
  assign new_n11637_ = new_n3794_ & new_n11614_;
  assign new_n11638_ = new_n11636_ & ~new_n11637_;
  assign new_n11639_ = ~new_n11624_ & ~new_n11625_;
  assign new_n11640_ = new_n11632_ & new_n11639_;
  assign new_n11641_ = new_n11638_ & new_n11640_;
  assign new_n11642_ = new_n4041_ & new_n11615_;
  assign new_n11643_ = new_n11641_ & ~new_n11642_;
  assign new_n11644_ = new_n3786_ & new_n11615_;
  assign new_n11645_ = lo0096 & new_n5140_;
  assign new_n11646_ = new_n11643_ & ~new_n11644_;
  assign new_n11647_ = ~new_n11645_ & new_n11646_;
  assign new_n11648_ = ~lo1044 & new_n11614_;
  assign new_n11649_ = new_n4007_ & new_n11648_;
  assign new_n11650_ = new_n3969_ & new_n11633_;
  assign new_n11651_ = ~new_n11649_ & ~new_n11650_;
  assign new_n11652_ = new_n3948_ & new_n11615_;
  assign new_n11653_ = lo0096 & ~new_n5216_;
  assign new_n11654_ = lo0096 & ~new_n4053_;
  assign new_n11655_ = ~li0583 & new_n11654_;
  assign new_n11656_ = lo0479 & new_n11655_;
  assign new_n11657_ = lo0096 & li0583;
  assign new_n11658_ = ~new_n11656_ & ~new_n11657_;
  assign new_n11659_ = new_n9406_ & ~new_n11658_;
  assign new_n11660_ = new_n4133_ & new_n11615_;
  assign new_n11661_ = ~new_n11659_ & ~new_n11660_;
  assign new_n11662_ = new_n11651_ & ~new_n11652_;
  assign new_n11663_ = ~new_n11653_ & new_n11662_;
  assign new_n11664_ = new_n11661_ & new_n11663_;
  assign new_n11665_ = new_n11647_ & new_n11664_;
  assign new_n11666_ = lo0096 & ~new_n5134_;
  assign new_n11667_ = ~new_n5201_ & new_n11633_;
  assign new_n11668_ = lo0096 & new_n5194_;
  assign new_n11669_ = ~new_n11615_ & ~new_n11668_;
  assign new_n11670_ = new_n3936_ & ~new_n11669_;
  assign new_n11671_ = new_n3625_ & new_n11615_;
  assign new_n11672_ = ~new_n11670_ & ~new_n11671_;
  assign new_n11673_ = lo0096 & new_n5818_;
  assign new_n11674_ = ~new_n5184_ & new_n11673_;
  assign new_n11675_ = lo0096 & new_n3706_;
  assign new_n11676_ = ~new_n11667_ & new_n11672_;
  assign new_n11677_ = ~new_n11674_ & new_n11676_;
  assign new_n11678_ = ~new_n11675_ & new_n11677_;
  assign new_n11679_ = new_n5133_ & new_n11666_;
  assign new_n11680_ = new_n11678_ & ~new_n11679_;
  assign new_n11681_ = lo0096 & new_n5505_;
  assign new_n11682_ = new_n11623_ & new_n11665_;
  assign new_n11683_ = new_n11680_ & new_n11682_;
  assign new_n11684_ = ~new_n11681_ & new_n11683_;
  assign new_n11685_ = new_n3804_ & new_n11615_;
  assign new_n11686_ = new_n3834_ & new_n11657_;
  assign new_n11687_ = new_n3678_ & new_n11686_;
  assign new_n11688_ = lo0096 & new_n5112_;
  assign new_n11689_ = new_n3810_ & new_n11633_;
  assign new_n11690_ = ~new_n11685_ & ~new_n11687_;
  assign new_n11691_ = ~new_n11688_ & new_n11690_;
  assign new_n11692_ = ~new_n11689_ & new_n11691_;
  assign new_n11693_ = ~new_n5105_ & new_n11633_;
  assign new_n11694_ = new_n11692_ & ~new_n11693_;
  assign new_n11695_ = new_n3815_ & new_n11614_;
  assign new_n11696_ = new_n4088_ & new_n11615_;
  assign new_n11697_ = ~new_n11695_ & ~new_n11696_;
  assign new_n11698_ = new_n3820_ & new_n11633_;
  assign new_n11699_ = new_n3870_ & new_n11648_;
  assign new_n11700_ = ~new_n11698_ & ~new_n11699_;
  assign new_n11701_ = ~new_n4069_ & new_n11615_;
  assign new_n11702_ = new_n11694_ & new_n11697_;
  assign new_n11703_ = new_n11700_ & new_n11702_;
  assign new_n11704_ = ~new_n11701_ & new_n11703_;
  assign new_n11705_ = ~new_n5096_ & new_n11633_;
  assign new_n11706_ = new_n3746_ & new_n11614_;
  assign new_n11707_ = ~new_n11705_ & ~new_n11706_;
  assign new_n11708_ = new_n4096_ & ~new_n11615_;
  assign new_n11709_ = ~lo0096 & ~new_n4096_;
  assign new_n11710_ = ~new_n11708_ & ~new_n11709_;
  assign new_n11711_ = ~lo0024 & ~lo0096;
  assign new_n11712_ = new_n4020_ & ~new_n11711_;
  assign new_n11713_ = new_n5090_ & new_n11710_;
  assign new_n11714_ = ~new_n11712_ & ~new_n11713_;
  assign new_n11715_ = lo0096 & new_n5071_;
  assign new_n11716_ = lo0096 & new_n4219_;
  assign new_n11717_ = ~new_n5074_ & new_n11716_;
  assign new_n11718_ = ~new_n5076_ & new_n11657_;
  assign new_n11719_ = ~new_n11717_ & ~new_n11718_;
  assign new_n11720_ = new_n4475_ & ~new_n11719_;
  assign new_n11721_ = lo0096 & new_n5083_;
  assign new_n11722_ = ~new_n11715_ & ~new_n11720_;
  assign new_n11723_ = ~new_n11721_ & new_n11722_;
  assign new_n11724_ = new_n5070_ & ~new_n11723_;
  assign new_n11725_ = new_n11704_ & new_n11707_;
  assign new_n11726_ = new_n11714_ & new_n11725_;
  assign new_n11727_ = ~new_n11724_ & new_n11726_;
  assign li0096 = ~new_n11684_ | ~new_n11727_;
  assign new_n11729_ = lo0097 & ~lo0314;
  assign new_n11730_ = ~lo0024 & lo0097;
  assign new_n11731_ = ~new_n5060_ & new_n11729_;
  assign new_n11732_ = new_n3940_ & new_n11730_;
  assign new_n11733_ = ~new_n11731_ & ~new_n11732_;
  assign new_n11734_ = lo0097 & ~lo0993;
  assign new_n11735_ = new_n3927_ & new_n11734_;
  assign new_n11736_ = new_n3953_ & new_n11730_;
  assign new_n11737_ = ~new_n11735_ & ~new_n11736_;
  assign new_n11738_ = new_n11733_ & new_n11737_;
  assign new_n11739_ = lo0097 & ~lo0841;
  assign new_n11740_ = new_n3763_ & new_n11739_;
  assign new_n11741_ = new_n3780_ & new_n11730_;
  assign new_n11742_ = ~new_n11740_ & ~new_n11741_;
  assign new_n11743_ = lo0097 & lo1076;
  assign new_n11744_ = new_n4050_ & new_n11730_;
  assign new_n11745_ = new_n3773_ & new_n11743_;
  assign new_n11746_ = ~new_n11744_ & ~new_n11745_;
  assign new_n11747_ = new_n3794_ & new_n11729_;
  assign new_n11748_ = ~new_n5460_ & new_n11729_;
  assign new_n11749_ = ~new_n11747_ & ~new_n11748_;
  assign new_n11750_ = new_n11746_ & new_n11749_;
  assign new_n11751_ = lo0097 & ~new_n4632_;
  assign new_n11752_ = lo0097 & new_n5155_;
  assign new_n11753_ = new_n3777_ & new_n11752_;
  assign new_n11754_ = new_n5565_ & new_n11751_;
  assign new_n11755_ = ~new_n11753_ & ~new_n11754_;
  assign new_n11756_ = new_n11742_ & new_n11750_;
  assign new_n11757_ = new_n11755_ & new_n11756_;
  assign new_n11758_ = new_n4041_ & new_n11730_;
  assign new_n11759_ = new_n11757_ & ~new_n11758_;
  assign new_n11760_ = new_n3786_ & new_n11730_;
  assign new_n11761_ = lo0097 & new_n5140_;
  assign new_n11762_ = new_n11759_ & ~new_n11760_;
  assign new_n11763_ = ~new_n11761_ & new_n11762_;
  assign new_n11764_ = ~lo1044 & new_n11729_;
  assign new_n11765_ = new_n4007_ & new_n11764_;
  assign new_n11766_ = new_n3969_ & new_n11739_;
  assign new_n11767_ = ~new_n11765_ & ~new_n11766_;
  assign new_n11768_ = new_n3948_ & new_n11730_;
  assign new_n11769_ = lo0097 & li0583;
  assign new_n11770_ = new_n3974_ & new_n11769_;
  assign new_n11771_ = ~new_n4135_ & new_n11770_;
  assign new_n11772_ = lo0097 & new_n5225_;
  assign new_n11773_ = ~new_n11771_ & ~new_n11772_;
  assign new_n11774_ = lo0097 & ~new_n5216_;
  assign new_n11775_ = new_n4133_ & new_n11730_;
  assign new_n11776_ = ~new_n11774_ & ~new_n11775_;
  assign new_n11777_ = new_n11767_ & ~new_n11768_;
  assign new_n11778_ = new_n11773_ & new_n11777_;
  assign new_n11779_ = new_n11776_ & new_n11778_;
  assign new_n11780_ = new_n11763_ & new_n11779_;
  assign new_n11781_ = lo0097 & ~new_n5134_;
  assign new_n11782_ = ~new_n5201_ & new_n11739_;
  assign new_n11783_ = lo0097 & new_n5194_;
  assign new_n11784_ = ~new_n11730_ & ~new_n11783_;
  assign new_n11785_ = new_n3936_ & ~new_n11784_;
  assign new_n11786_ = new_n3625_ & new_n11730_;
  assign new_n11787_ = ~new_n11785_ & ~new_n11786_;
  assign new_n11788_ = lo0097 & new_n5818_;
  assign new_n11789_ = ~new_n5184_ & new_n11788_;
  assign new_n11790_ = lo0097 & new_n3706_;
  assign new_n11791_ = ~new_n11782_ & new_n11787_;
  assign new_n11792_ = ~new_n11789_ & new_n11791_;
  assign new_n11793_ = ~new_n11790_ & new_n11792_;
  assign new_n11794_ = new_n5133_ & new_n11781_;
  assign new_n11795_ = new_n11793_ & ~new_n11794_;
  assign new_n11796_ = lo0097 & new_n5505_;
  assign new_n11797_ = new_n11738_ & new_n11780_;
  assign new_n11798_ = new_n11795_ & new_n11797_;
  assign new_n11799_ = ~new_n11796_ & new_n11798_;
  assign new_n11800_ = new_n3804_ & new_n11730_;
  assign new_n11801_ = new_n3834_ & new_n11769_;
  assign new_n11802_ = new_n3678_ & new_n11801_;
  assign new_n11803_ = lo0097 & new_n5112_;
  assign new_n11804_ = new_n3810_ & new_n11739_;
  assign new_n11805_ = ~new_n11800_ & ~new_n11802_;
  assign new_n11806_ = ~new_n11803_ & new_n11805_;
  assign new_n11807_ = ~new_n11804_ & new_n11806_;
  assign new_n11808_ = ~new_n5105_ & new_n11739_;
  assign new_n11809_ = new_n11807_ & ~new_n11808_;
  assign new_n11810_ = new_n3815_ & new_n11729_;
  assign new_n11811_ = new_n4088_ & new_n11730_;
  assign new_n11812_ = ~new_n11810_ & ~new_n11811_;
  assign new_n11813_ = new_n3820_ & new_n11739_;
  assign new_n11814_ = new_n3870_ & new_n11764_;
  assign new_n11815_ = ~new_n11813_ & ~new_n11814_;
  assign new_n11816_ = ~new_n4069_ & new_n11730_;
  assign new_n11817_ = new_n11809_ & new_n11812_;
  assign new_n11818_ = new_n11815_ & new_n11817_;
  assign new_n11819_ = ~new_n11816_ & new_n11818_;
  assign new_n11820_ = new_n4020_ & new_n11730_;
  assign new_n11821_ = ~new_n5096_ & new_n11739_;
  assign new_n11822_ = ~new_n11820_ & ~new_n11821_;
  assign new_n11823_ = ~new_n4096_ & new_n11730_;
  assign new_n11824_ = lo0097 & ~new_n11730_;
  assign new_n11825_ = ~new_n11823_ & ~new_n11824_;
  assign new_n11826_ = new_n5090_ & ~new_n11825_;
  assign new_n11827_ = new_n3746_ & new_n11729_;
  assign new_n11828_ = ~new_n11826_ & ~new_n11827_;
  assign new_n11829_ = lo0097 & new_n5071_;
  assign new_n11830_ = lo0097 & ~new_n5074_;
  assign new_n11831_ = new_n5074_ & new_n8961_;
  assign new_n11832_ = ~new_n11830_ & ~new_n11831_;
  assign new_n11833_ = ~new_n5076_ & new_n11769_;
  assign new_n11834_ = new_n4219_ & ~new_n11832_;
  assign new_n11835_ = ~new_n11833_ & ~new_n11834_;
  assign new_n11836_ = new_n4475_ & ~new_n11835_;
  assign new_n11837_ = lo0097 & new_n5083_;
  assign new_n11838_ = ~new_n11829_ & ~new_n11836_;
  assign new_n11839_ = ~new_n11837_ & new_n11838_;
  assign new_n11840_ = new_n5070_ & ~new_n11839_;
  assign new_n11841_ = new_n11819_ & new_n11822_;
  assign new_n11842_ = new_n11828_ & new_n11841_;
  assign new_n11843_ = ~new_n11840_ & new_n11842_;
  assign li0097 = ~new_n11799_ | ~new_n11843_;
  assign new_n11845_ = lo0098 & new_n4001_;
  assign new_n11846_ = lo0098 & ~lo0841;
  assign new_n11847_ = ~new_n5201_ & new_n11846_;
  assign new_n11848_ = ~lo0024 & lo0098;
  assign new_n11849_ = lo0098 & new_n5194_;
  assign new_n11850_ = ~new_n11848_ & ~new_n11849_;
  assign new_n11851_ = new_n3936_ & ~new_n11850_;
  assign new_n11852_ = new_n3625_ & new_n11848_;
  assign new_n11853_ = ~new_n11851_ & ~new_n11852_;
  assign new_n11854_ = ~new_n11847_ & new_n11853_;
  assign new_n11855_ = new_n5230_ & new_n11845_;
  assign new_n11856_ = new_n11854_ & ~new_n11855_;
  assign new_n11857_ = new_n3763_ & new_n11846_;
  assign new_n11858_ = new_n3780_ & new_n11848_;
  assign new_n11859_ = ~new_n11857_ & ~new_n11858_;
  assign new_n11860_ = lo0098 & lo1076;
  assign new_n11861_ = new_n4050_ & new_n11848_;
  assign new_n11862_ = new_n3773_ & new_n11860_;
  assign new_n11863_ = ~new_n11861_ & ~new_n11862_;
  assign new_n11864_ = lo0098 & ~lo0314;
  assign new_n11865_ = new_n3794_ & new_n11864_;
  assign new_n11866_ = ~new_n5460_ & new_n11864_;
  assign new_n11867_ = ~new_n11865_ & ~new_n11866_;
  assign new_n11868_ = new_n11863_ & new_n11867_;
  assign new_n11869_ = lo0098 & ~new_n4632_;
  assign new_n11870_ = lo0098 & new_n5155_;
  assign new_n11871_ = new_n3777_ & new_n11870_;
  assign new_n11872_ = new_n5565_ & new_n11869_;
  assign new_n11873_ = ~new_n11871_ & ~new_n11872_;
  assign new_n11874_ = new_n11859_ & new_n11868_;
  assign new_n11875_ = new_n11873_ & new_n11874_;
  assign new_n11876_ = new_n4041_ & new_n11848_;
  assign new_n11877_ = new_n11875_ & ~new_n11876_;
  assign new_n11878_ = new_n3786_ & new_n11848_;
  assign new_n11879_ = lo0098 & new_n5140_;
  assign new_n11880_ = new_n11877_ & ~new_n11878_;
  assign new_n11881_ = ~new_n11879_ & new_n11880_;
  assign new_n11882_ = new_n3969_ & new_n11846_;
  assign new_n11883_ = new_n3948_ & new_n11848_;
  assign new_n11884_ = ~new_n11882_ & ~new_n11883_;
  assign new_n11885_ = new_n4133_ & new_n11848_;
  assign new_n11886_ = lo0098 & li0583;
  assign new_n11887_ = new_n3974_ & new_n11886_;
  assign new_n11888_ = ~new_n4135_ & new_n11887_;
  assign new_n11889_ = lo0098 & new_n5225_;
  assign new_n11890_ = ~new_n11888_ & ~new_n11889_;
  assign new_n11891_ = ~lo0098 & ~lo0314;
  assign new_n11892_ = ~lo1044 & ~new_n11891_;
  assign new_n11893_ = new_n4007_ & new_n11892_;
  assign new_n11894_ = lo0098 & ~new_n5216_;
  assign new_n11895_ = ~new_n11893_ & ~new_n11894_;
  assign new_n11896_ = new_n11884_ & ~new_n11885_;
  assign new_n11897_ = new_n11890_ & new_n11896_;
  assign new_n11898_ = new_n11895_ & new_n11897_;
  assign new_n11899_ = new_n11881_ & new_n11898_;
  assign new_n11900_ = lo0098 & new_n5608_;
  assign new_n11901_ = ~new_n5184_ & new_n11900_;
  assign new_n11902_ = lo0098 & new_n3706_;
  assign new_n11903_ = lo0098 & new_n5133_;
  assign new_n11904_ = ~new_n5134_ & new_n11903_;
  assign new_n11905_ = ~new_n11901_ & ~new_n11902_;
  assign new_n11906_ = ~new_n11904_ & new_n11905_;
  assign new_n11907_ = ~new_n5060_ & new_n11864_;
  assign new_n11908_ = new_n3940_ & new_n11848_;
  assign new_n11909_ = ~new_n11907_ & ~new_n11908_;
  assign new_n11910_ = lo0098 & ~lo0993;
  assign new_n11911_ = new_n3927_ & new_n11910_;
  assign new_n11912_ = new_n3953_ & new_n11848_;
  assign new_n11913_ = ~new_n11911_ & ~new_n11912_;
  assign new_n11914_ = new_n11909_ & new_n11913_;
  assign new_n11915_ = new_n11856_ & new_n11899_;
  assign new_n11916_ = new_n11906_ & new_n11915_;
  assign new_n11917_ = new_n11914_ & new_n11916_;
  assign new_n11918_ = ~new_n5096_ & new_n11846_;
  assign new_n11919_ = new_n4020_ & new_n11848_;
  assign new_n11920_ = ~new_n11918_ & ~new_n11919_;
  assign new_n11921_ = lo0098 & new_n5071_;
  assign new_n11922_ = lo0098 & lo0786;
  assign new_n11923_ = ~new_n5076_ & new_n11886_;
  assign new_n11924_ = lo0098 & new_n5545_;
  assign new_n11925_ = ~new_n11923_ & ~new_n11924_;
  assign new_n11926_ = new_n4475_ & ~new_n11925_;
  assign new_n11927_ = new_n5082_ & new_n11922_;
  assign new_n11928_ = ~new_n11926_ & ~new_n11927_;
  assign new_n11929_ = ~new_n11921_ & new_n11928_;
  assign new_n11930_ = new_n5070_ & ~new_n11929_;
  assign new_n11931_ = new_n3746_ & new_n11864_;
  assign new_n11932_ = ~new_n4096_ & new_n11848_;
  assign new_n11933_ = lo0098 & ~new_n11848_;
  assign new_n11934_ = ~new_n11932_ & ~new_n11933_;
  assign new_n11935_ = new_n5090_ & ~new_n11934_;
  assign new_n11936_ = ~new_n11931_ & ~new_n11935_;
  assign new_n11937_ = ~new_n11930_ & new_n11936_;
  assign new_n11938_ = new_n11920_ & new_n11937_;
  assign new_n11939_ = new_n3870_ & new_n11892_;
  assign new_n11940_ = new_n3834_ & new_n11886_;
  assign new_n11941_ = new_n3678_ & new_n11940_;
  assign new_n11942_ = lo0098 & new_n5112_;
  assign new_n11943_ = new_n3810_ & new_n11846_;
  assign new_n11944_ = ~new_n11939_ & ~new_n11941_;
  assign new_n11945_ = ~new_n11942_ & new_n11944_;
  assign new_n11946_ = ~new_n11943_ & new_n11945_;
  assign new_n11947_ = ~new_n5105_ & new_n11846_;
  assign new_n11948_ = new_n11946_ & ~new_n11947_;
  assign new_n11949_ = new_n3815_ & new_n11864_;
  assign new_n11950_ = new_n4088_ & new_n11848_;
  assign new_n11951_ = ~new_n11949_ & ~new_n11950_;
  assign new_n11952_ = new_n3820_ & new_n11846_;
  assign new_n11953_ = new_n3618_ & new_n11848_;
  assign new_n11954_ = ~new_n11952_ & ~new_n11953_;
  assign new_n11955_ = ~new_n5394_ & new_n11848_;
  assign new_n11956_ = new_n11954_ & ~new_n11955_;
  assign new_n11957_ = new_n11938_ & new_n11948_;
  assign new_n11958_ = new_n11951_ & new_n11957_;
  assign new_n11959_ = new_n11956_ & new_n11958_;
  assign li0098 = ~new_n11917_ | ~new_n11959_;
  assign new_n11961_ = lo0099 & ~new_n6030_;
  assign new_n11962_ = ~new_n6044_ & ~new_n11961_;
  assign new_n11963_ = new_n6028_ & ~new_n11962_;
  assign new_n11964_ = lo0099 & ~new_n6028_;
  assign new_n11965_ = ~new_n11963_ & ~new_n11964_;
  assign new_n11966_ = ~lo0039 & ~lo0072;
  assign new_n11967_ = ~lo0072 & ~new_n5253_;
  assign new_n11968_ = lo0039 & new_n11967_;
  assign new_n11969_ = ~new_n11965_ & new_n11966_;
  assign new_n11970_ = new_n6038_ & new_n11968_;
  assign li0099 = new_n11969_ | new_n11970_;
  assign new_n11972_ = lo0100 & ~lo0314;
  assign new_n11973_ = ~lo0024 & lo0100;
  assign new_n11974_ = ~new_n5060_ & new_n11972_;
  assign new_n11975_ = new_n3940_ & new_n11973_;
  assign new_n11976_ = ~new_n11974_ & ~new_n11975_;
  assign new_n11977_ = lo0100 & ~lo0993;
  assign new_n11978_ = new_n3927_ & new_n11977_;
  assign new_n11979_ = new_n3953_ & new_n11973_;
  assign new_n11980_ = ~new_n11978_ & ~new_n11979_;
  assign new_n11981_ = lo0100 & new_n5071_;
  assign new_n11982_ = lo0100 & new_n4219_;
  assign new_n11983_ = lo0100 & li0583;
  assign new_n11984_ = ~new_n5074_ & new_n11982_;
  assign new_n11985_ = ~new_n5076_ & new_n11983_;
  assign new_n11986_ = ~new_n11984_ & ~new_n11985_;
  assign new_n11987_ = new_n4475_ & ~new_n11986_;
  assign new_n11988_ = lo0100 & new_n5083_;
  assign new_n11989_ = ~new_n11981_ & ~new_n11987_;
  assign new_n11990_ = ~new_n11988_ & new_n11989_;
  assign new_n11991_ = new_n3746_ & new_n11972_;
  assign new_n11992_ = ~new_n4096_ & new_n11973_;
  assign new_n11993_ = lo0100 & ~new_n11973_;
  assign new_n11994_ = ~new_n11992_ & ~new_n11993_;
  assign new_n11995_ = new_n5090_ & ~new_n11994_;
  assign new_n11996_ = ~new_n11991_ & ~new_n11995_;
  assign new_n11997_ = new_n5070_ & ~new_n11990_;
  assign new_n11998_ = new_n11996_ & ~new_n11997_;
  assign new_n11999_ = lo0100 & ~lo0841;
  assign new_n12000_ = new_n4020_ & new_n11973_;
  assign new_n12001_ = ~new_n5096_ & new_n11999_;
  assign new_n12002_ = ~new_n12000_ & ~new_n12001_;
  assign new_n12003_ = new_n11976_ & new_n11980_;
  assign new_n12004_ = new_n11998_ & new_n12003_;
  assign new_n12005_ = new_n12002_ & new_n12004_;
  assign new_n12006_ = new_n3804_ & new_n11973_;
  assign new_n12007_ = new_n3834_ & new_n11983_;
  assign new_n12008_ = new_n3678_ & new_n12007_;
  assign new_n12009_ = lo0100 & new_n5112_;
  assign new_n12010_ = new_n3810_ & new_n11999_;
  assign new_n12011_ = ~new_n12006_ & ~new_n12008_;
  assign new_n12012_ = ~new_n12009_ & new_n12011_;
  assign new_n12013_ = ~new_n12010_ & new_n12012_;
  assign new_n12014_ = ~new_n5105_ & new_n11999_;
  assign new_n12015_ = new_n12013_ & ~new_n12014_;
  assign new_n12016_ = new_n3815_ & new_n11972_;
  assign new_n12017_ = new_n4088_ & new_n11973_;
  assign new_n12018_ = ~new_n12016_ & ~new_n12017_;
  assign new_n12019_ = ~lo1044 & new_n11972_;
  assign new_n12020_ = new_n3820_ & new_n11999_;
  assign new_n12021_ = new_n3870_ & new_n12019_;
  assign new_n12022_ = ~new_n12020_ & ~new_n12021_;
  assign new_n12023_ = ~new_n4069_ & new_n11973_;
  assign new_n12024_ = new_n12015_ & new_n12018_;
  assign new_n12025_ = new_n12022_ & new_n12024_;
  assign new_n12026_ = ~new_n12023_ & new_n12025_;
  assign new_n12027_ = lo0100 & new_n5135_;
  assign new_n12028_ = lo0100 & lo1076;
  assign new_n12029_ = lo0024 & ~new_n5169_;
  assign new_n12030_ = li0683 & new_n12029_;
  assign new_n12031_ = ~new_n11973_ & ~new_n12030_;
  assign new_n12032_ = new_n4050_ & ~new_n12031_;
  assign new_n12033_ = new_n3773_ & new_n12028_;
  assign new_n12034_ = ~new_n12032_ & ~new_n12033_;
  assign new_n12035_ = lo0100 & new_n5155_;
  assign new_n12036_ = new_n3777_ & new_n12035_;
  assign new_n12037_ = lo0100 & ~new_n4632_;
  assign new_n12038_ = new_n5565_ & new_n12037_;
  assign new_n12039_ = ~new_n12036_ & ~new_n12038_;
  assign new_n12040_ = ~new_n5460_ & new_n11972_;
  assign new_n12041_ = new_n12039_ & ~new_n12040_;
  assign new_n12042_ = new_n3780_ & new_n11973_;
  assign new_n12043_ = new_n3763_ & new_n11999_;
  assign new_n12044_ = ~new_n12042_ & ~new_n12043_;
  assign new_n12045_ = new_n3794_ & new_n11972_;
  assign new_n12046_ = new_n12034_ & new_n12041_;
  assign new_n12047_ = new_n12044_ & new_n12046_;
  assign new_n12048_ = ~new_n12045_ & new_n12047_;
  assign new_n12049_ = new_n4041_ & new_n11973_;
  assign new_n12050_ = new_n12048_ & ~new_n12049_;
  assign new_n12051_ = lo0100 & new_n5140_;
  assign new_n12052_ = new_n3786_ & new_n11973_;
  assign new_n12053_ = ~new_n12027_ & new_n12050_;
  assign new_n12054_ = ~new_n12051_ & new_n12053_;
  assign new_n12055_ = ~new_n12052_ & new_n12054_;
  assign new_n12056_ = lo0100 & new_n5194_;
  assign new_n12057_ = ~new_n11973_ & ~new_n12056_;
  assign new_n12058_ = new_n3936_ & ~new_n12057_;
  assign new_n12059_ = new_n3625_ & new_n11973_;
  assign new_n12060_ = ~new_n12058_ & ~new_n12059_;
  assign new_n12061_ = lo0100 & new_n3706_;
  assign new_n12062_ = lo0100 & new_n5608_;
  assign new_n12063_ = ~new_n5184_ & new_n12062_;
  assign new_n12064_ = new_n12060_ & ~new_n12061_;
  assign new_n12065_ = ~new_n12063_ & new_n12064_;
  assign new_n12066_ = ~new_n5201_ & new_n11999_;
  assign new_n12067_ = new_n12065_ & ~new_n12066_;
  assign new_n12068_ = lo0100 & new_n5505_;
  assign new_n12069_ = new_n4007_ & new_n12019_;
  assign new_n12070_ = new_n3969_ & new_n11999_;
  assign new_n12071_ = ~new_n12069_ & ~new_n12070_;
  assign new_n12072_ = lo0100 & ~new_n5216_;
  assign new_n12073_ = new_n4133_ & new_n11973_;
  assign new_n12074_ = ~new_n12072_ & ~new_n12073_;
  assign new_n12075_ = new_n3974_ & new_n11983_;
  assign new_n12076_ = ~new_n4135_ & new_n12075_;
  assign new_n12077_ = lo0100 & new_n5225_;
  assign new_n12078_ = new_n12074_ & ~new_n12076_;
  assign new_n12079_ = ~new_n12077_ & new_n12078_;
  assign new_n12080_ = new_n3948_ & new_n11973_;
  assign new_n12081_ = new_n12079_ & ~new_n12080_;
  assign new_n12082_ = new_n12067_ & ~new_n12068_;
  assign new_n12083_ = new_n12071_ & new_n12082_;
  assign new_n12084_ = new_n12081_ & new_n12083_;
  assign new_n12085_ = new_n12005_ & new_n12026_;
  assign new_n12086_ = new_n12055_ & new_n12085_;
  assign li0100 = ~new_n12084_ | ~new_n12086_;
  assign new_n12088_ = lo0044 & lo0101;
  assign new_n12089_ = ~new_n6029_ & ~new_n12088_;
  assign new_n12090_ = new_n6028_ & ~new_n12089_;
  assign new_n12091_ = lo0101 & ~new_n6028_;
  assign new_n12092_ = ~new_n12090_ & ~new_n12091_;
  assign new_n12093_ = new_n11966_ & ~new_n12092_;
  assign new_n12094_ = new_n6102_ & new_n11968_;
  assign li0101 = new_n12093_ | new_n12094_;
  assign new_n12096_ = lo0102 & ~lo0841;
  assign new_n12097_ = lo0102 & new_n5818_;
  assign new_n12098_ = ~new_n5184_ & new_n12097_;
  assign new_n12099_ = lo0102 & new_n3706_;
  assign new_n12100_ = ~lo0024 & lo0102;
  assign new_n12101_ = lo0102 & new_n5194_;
  assign new_n12102_ = ~new_n12100_ & ~new_n12101_;
  assign new_n12103_ = new_n3936_ & ~new_n12102_;
  assign new_n12104_ = new_n3625_ & new_n12100_;
  assign new_n12105_ = ~new_n12103_ & ~new_n12104_;
  assign new_n12106_ = ~new_n12098_ & ~new_n12099_;
  assign new_n12107_ = new_n12105_ & new_n12106_;
  assign new_n12108_ = ~new_n5201_ & new_n12096_;
  assign new_n12109_ = new_n12107_ & ~new_n12108_;
  assign new_n12110_ = lo0102 & ~lo0993;
  assign new_n12111_ = new_n3927_ & new_n12110_;
  assign new_n12112_ = new_n3953_ & new_n12100_;
  assign new_n12113_ = ~new_n12111_ & ~new_n12112_;
  assign new_n12114_ = new_n12109_ & new_n12113_;
  assign new_n12115_ = new_n3804_ & new_n12100_;
  assign new_n12116_ = lo0102 & li0583;
  assign new_n12117_ = new_n3834_ & new_n12116_;
  assign new_n12118_ = new_n3678_ & new_n12117_;
  assign new_n12119_ = lo0102 & new_n5112_;
  assign new_n12120_ = new_n3810_ & new_n12096_;
  assign new_n12121_ = ~new_n12115_ & ~new_n12118_;
  assign new_n12122_ = ~new_n12119_ & new_n12121_;
  assign new_n12123_ = ~new_n12120_ & new_n12122_;
  assign new_n12124_ = ~new_n5105_ & new_n12096_;
  assign new_n12125_ = new_n12123_ & ~new_n12124_;
  assign new_n12126_ = new_n4050_ & new_n12100_;
  assign new_n12127_ = lo0102 & new_n5562_;
  assign new_n12128_ = lo0102 & ~lo0314;
  assign new_n12129_ = lo0102 & new_n5155_;
  assign new_n12130_ = new_n3777_ & new_n12129_;
  assign new_n12131_ = lo0102 & ~new_n4632_;
  assign new_n12132_ = new_n5565_ & new_n12131_;
  assign new_n12133_ = ~new_n12130_ & ~new_n12132_;
  assign new_n12134_ = ~new_n5460_ & new_n12128_;
  assign new_n12135_ = new_n12133_ & ~new_n12134_;
  assign new_n12136_ = new_n3763_ & new_n12096_;
  assign new_n12137_ = new_n3780_ & new_n12100_;
  assign new_n12138_ = ~new_n12136_ & ~new_n12137_;
  assign new_n12139_ = new_n3794_ & new_n12128_;
  assign new_n12140_ = new_n12138_ & ~new_n12139_;
  assign new_n12141_ = ~new_n12126_ & ~new_n12127_;
  assign new_n12142_ = new_n12135_ & new_n12141_;
  assign new_n12143_ = new_n12140_ & new_n12142_;
  assign new_n12144_ = new_n4041_ & new_n12100_;
  assign new_n12145_ = new_n12143_ & ~new_n12144_;
  assign new_n12146_ = new_n3815_ & new_n12128_;
  assign new_n12147_ = new_n4088_ & new_n12100_;
  assign new_n12148_ = ~new_n12146_ & ~new_n12147_;
  assign new_n12149_ = lo0102 & new_n3678_;
  assign new_n12150_ = new_n3786_ & new_n12100_;
  assign new_n12151_ = new_n5139_ & new_n12149_;
  assign new_n12152_ = ~new_n12150_ & ~new_n12151_;
  assign new_n12153_ = new_n12125_ & new_n12145_;
  assign new_n12154_ = new_n12148_ & new_n12153_;
  assign new_n12155_ = new_n12152_ & new_n12154_;
  assign new_n12156_ = new_n12114_ & new_n12155_;
  assign new_n12157_ = new_n4020_ & new_n12100_;
  assign new_n12158_ = ~lo1044 & new_n12128_;
  assign new_n12159_ = new_n3820_ & new_n12096_;
  assign new_n12160_ = new_n3870_ & new_n12158_;
  assign new_n12161_ = ~new_n12159_ & ~new_n12160_;
  assign new_n12162_ = ~new_n4069_ & new_n12100_;
  assign new_n12163_ = ~new_n5096_ & new_n12096_;
  assign new_n12164_ = ~new_n12157_ & new_n12161_;
  assign new_n12165_ = ~new_n12162_ & new_n12164_;
  assign new_n12166_ = ~new_n12163_ & new_n12165_;
  assign new_n12167_ = new_n3746_ & new_n12128_;
  assign new_n12168_ = ~new_n4096_ & new_n12100_;
  assign new_n12169_ = lo0102 & ~new_n12100_;
  assign new_n12170_ = ~new_n12168_ & ~new_n12169_;
  assign new_n12171_ = new_n5090_ & ~new_n12170_;
  assign new_n12172_ = ~new_n12167_ & ~new_n12171_;
  assign new_n12173_ = new_n12166_ & new_n12172_;
  assign new_n12174_ = lo0102 & new_n5505_;
  assign new_n12175_ = new_n12173_ & ~new_n12174_;
  assign new_n12176_ = lo0102 & ~new_n5216_;
  assign new_n12177_ = new_n4133_ & new_n12100_;
  assign new_n12178_ = ~new_n12176_ & ~new_n12177_;
  assign new_n12179_ = new_n3974_ & new_n12116_;
  assign new_n12180_ = ~new_n4135_ & new_n12179_;
  assign new_n12181_ = lo0102 & new_n5225_;
  assign new_n12182_ = new_n12178_ & ~new_n12180_;
  assign new_n12183_ = ~new_n12181_ & new_n12182_;
  assign new_n12184_ = new_n3948_ & new_n12100_;
  assign new_n12185_ = new_n12183_ & ~new_n12184_;
  assign new_n12186_ = new_n4007_ & new_n12158_;
  assign new_n12187_ = new_n3969_ & new_n12096_;
  assign new_n12188_ = ~new_n12186_ & ~new_n12187_;
  assign new_n12189_ = ~new_n3922_ & new_n12185_;
  assign new_n12190_ = new_n12188_ & new_n12189_;
  assign new_n12191_ = lo0102 & new_n5071_;
  assign new_n12192_ = lo0102 & new_n4219_;
  assign new_n12193_ = ~new_n5074_ & new_n12192_;
  assign new_n12194_ = ~new_n5076_ & new_n12116_;
  assign new_n12195_ = ~new_n12193_ & ~new_n12194_;
  assign new_n12196_ = new_n4475_ & ~new_n12195_;
  assign new_n12197_ = lo0102 & new_n5083_;
  assign new_n12198_ = ~new_n12191_ & ~new_n12196_;
  assign new_n12199_ = ~new_n12197_ & new_n12198_;
  assign new_n12200_ = new_n5070_ & ~new_n12199_;
  assign new_n12201_ = new_n12190_ & ~new_n12200_;
  assign new_n12202_ = lo0102 & new_n5135_;
  assign new_n12203_ = new_n3940_ & new_n12100_;
  assign new_n12204_ = ~new_n12202_ & ~new_n12203_;
  assign new_n12205_ = ~new_n5060_ & new_n12128_;
  assign new_n12206_ = new_n12204_ & ~new_n12205_;
  assign new_n12207_ = new_n12156_ & new_n12175_;
  assign new_n12208_ = new_n12201_ & new_n12207_;
  assign li0102 = ~new_n12206_ | ~new_n12208_;
  assign new_n12210_ = lo0103 & ~lo0841;
  assign new_n12211_ = lo0103 & new_n5818_;
  assign new_n12212_ = ~new_n5184_ & new_n12211_;
  assign new_n12213_ = lo0103 & new_n3706_;
  assign new_n12214_ = ~lo0024 & lo0103;
  assign new_n12215_ = lo0103 & new_n5194_;
  assign new_n12216_ = ~new_n12214_ & ~new_n12215_;
  assign new_n12217_ = new_n3936_ & ~new_n12216_;
  assign new_n12218_ = new_n3625_ & new_n12214_;
  assign new_n12219_ = ~new_n12217_ & ~new_n12218_;
  assign new_n12220_ = ~new_n12212_ & ~new_n12213_;
  assign new_n12221_ = new_n12219_ & new_n12220_;
  assign new_n12222_ = ~new_n5201_ & new_n12210_;
  assign new_n12223_ = new_n12221_ & ~new_n12222_;
  assign new_n12224_ = lo0103 & ~lo0993;
  assign new_n12225_ = new_n3927_ & new_n12224_;
  assign new_n12226_ = new_n3953_ & new_n12214_;
  assign new_n12227_ = ~new_n12225_ & ~new_n12226_;
  assign new_n12228_ = new_n12223_ & new_n12227_;
  assign new_n12229_ = new_n3804_ & new_n12214_;
  assign new_n12230_ = lo0103 & li0583;
  assign new_n12231_ = new_n3834_ & new_n12230_;
  assign new_n12232_ = new_n3678_ & new_n12231_;
  assign new_n12233_ = lo0103 & new_n5112_;
  assign new_n12234_ = new_n3810_ & new_n12210_;
  assign new_n12235_ = ~new_n12229_ & ~new_n12232_;
  assign new_n12236_ = ~new_n12233_ & new_n12235_;
  assign new_n12237_ = ~new_n12234_ & new_n12236_;
  assign new_n12238_ = ~new_n5105_ & new_n12210_;
  assign new_n12239_ = new_n12237_ & ~new_n12238_;
  assign new_n12240_ = new_n4050_ & new_n12214_;
  assign new_n12241_ = lo0103 & new_n5562_;
  assign new_n12242_ = lo0103 & ~lo0314;
  assign new_n12243_ = lo0103 & new_n5155_;
  assign new_n12244_ = new_n3777_ & new_n12243_;
  assign new_n12245_ = lo0103 & ~new_n4632_;
  assign new_n12246_ = new_n5565_ & new_n12245_;
  assign new_n12247_ = ~new_n12244_ & ~new_n12246_;
  assign new_n12248_ = ~new_n5460_ & new_n12242_;
  assign new_n12249_ = new_n12247_ & ~new_n12248_;
  assign new_n12250_ = new_n3763_ & new_n12210_;
  assign new_n12251_ = new_n3780_ & new_n12214_;
  assign new_n12252_ = ~new_n12250_ & ~new_n12251_;
  assign new_n12253_ = new_n3794_ & new_n12242_;
  assign new_n12254_ = new_n12252_ & ~new_n12253_;
  assign new_n12255_ = ~new_n12240_ & ~new_n12241_;
  assign new_n12256_ = new_n12249_ & new_n12255_;
  assign new_n12257_ = new_n12254_ & new_n12256_;
  assign new_n12258_ = new_n4041_ & new_n12214_;
  assign new_n12259_ = new_n12257_ & ~new_n12258_;
  assign new_n12260_ = new_n3815_ & new_n12242_;
  assign new_n12261_ = new_n4088_ & new_n12214_;
  assign new_n12262_ = ~new_n12260_ & ~new_n12261_;
  assign new_n12263_ = lo0103 & new_n3678_;
  assign new_n12264_ = new_n3786_ & new_n12214_;
  assign new_n12265_ = new_n5139_ & new_n12263_;
  assign new_n12266_ = ~new_n12264_ & ~new_n12265_;
  assign new_n12267_ = new_n12239_ & new_n12259_;
  assign new_n12268_ = new_n12262_ & new_n12267_;
  assign new_n12269_ = new_n12266_ & new_n12268_;
  assign new_n12270_ = new_n12228_ & new_n12269_;
  assign new_n12271_ = new_n4020_ & new_n12214_;
  assign new_n12272_ = ~lo1044 & new_n12242_;
  assign new_n12273_ = new_n3820_ & new_n12210_;
  assign new_n12274_ = new_n3870_ & new_n12272_;
  assign new_n12275_ = ~new_n12273_ & ~new_n12274_;
  assign new_n12276_ = ~new_n4069_ & new_n12214_;
  assign new_n12277_ = ~new_n5096_ & new_n12210_;
  assign new_n12278_ = ~new_n12271_ & new_n12275_;
  assign new_n12279_ = ~new_n12276_ & new_n12278_;
  assign new_n12280_ = ~new_n12277_ & new_n12279_;
  assign new_n12281_ = new_n3746_ & new_n12242_;
  assign new_n12282_ = ~new_n4096_ & new_n12214_;
  assign new_n12283_ = lo0103 & ~new_n12214_;
  assign new_n12284_ = ~new_n12282_ & ~new_n12283_;
  assign new_n12285_ = new_n5090_ & ~new_n12284_;
  assign new_n12286_ = ~new_n12281_ & ~new_n12285_;
  assign new_n12287_ = new_n12280_ & new_n12286_;
  assign new_n12288_ = lo0103 & new_n5505_;
  assign new_n12289_ = new_n12287_ & ~new_n12288_;
  assign new_n12290_ = lo0103 & ~new_n5216_;
  assign new_n12291_ = new_n4133_ & new_n12214_;
  assign new_n12292_ = ~new_n12290_ & ~new_n12291_;
  assign new_n12293_ = new_n3974_ & new_n12230_;
  assign new_n12294_ = ~new_n4135_ & new_n12293_;
  assign new_n12295_ = lo0103 & new_n5225_;
  assign new_n12296_ = new_n12292_ & ~new_n12294_;
  assign new_n12297_ = ~new_n12295_ & new_n12296_;
  assign new_n12298_ = new_n3948_ & new_n12214_;
  assign new_n12299_ = new_n12297_ & ~new_n12298_;
  assign new_n12300_ = new_n4007_ & new_n12272_;
  assign new_n12301_ = new_n3969_ & new_n12210_;
  assign new_n12302_ = ~new_n12300_ & ~new_n12301_;
  assign new_n12303_ = ~new_n3962_ & new_n12299_;
  assign new_n12304_ = new_n12302_ & new_n12303_;
  assign new_n12305_ = lo0103 & new_n5071_;
  assign new_n12306_ = lo0103 & new_n4219_;
  assign new_n12307_ = ~new_n5074_ & new_n12306_;
  assign new_n12308_ = ~new_n5076_ & new_n12230_;
  assign new_n12309_ = ~new_n12307_ & ~new_n12308_;
  assign new_n12310_ = new_n4475_ & ~new_n12309_;
  assign new_n12311_ = lo0103 & new_n5083_;
  assign new_n12312_ = ~new_n12305_ & ~new_n12310_;
  assign new_n12313_ = ~new_n12311_ & new_n12312_;
  assign new_n12314_ = new_n5070_ & ~new_n12313_;
  assign new_n12315_ = new_n12304_ & ~new_n12314_;
  assign new_n12316_ = lo0103 & new_n5135_;
  assign new_n12317_ = new_n3940_ & new_n12214_;
  assign new_n12318_ = ~new_n12316_ & ~new_n12317_;
  assign new_n12319_ = ~new_n5060_ & new_n12242_;
  assign new_n12320_ = new_n12318_ & ~new_n12319_;
  assign new_n12321_ = new_n12270_ & new_n12289_;
  assign new_n12322_ = new_n12315_ & new_n12321_;
  assign li0103 = ~new_n12320_ | ~new_n12322_;
  assign new_n12324_ = lo0104 & ~lo0314;
  assign new_n12325_ = ~lo0024 & lo0104;
  assign new_n12326_ = ~new_n5060_ & new_n12324_;
  assign new_n12327_ = new_n3940_ & new_n12325_;
  assign new_n12328_ = ~new_n12326_ & ~new_n12327_;
  assign new_n12329_ = lo0104 & ~lo0993;
  assign new_n12330_ = new_n3927_ & new_n12329_;
  assign new_n12331_ = new_n3953_ & new_n12325_;
  assign new_n12332_ = ~new_n12330_ & ~new_n12331_;
  assign new_n12333_ = lo0104 & new_n5071_;
  assign new_n12334_ = lo0104 & new_n4219_;
  assign new_n12335_ = lo0104 & li0583;
  assign new_n12336_ = ~new_n5074_ & new_n12334_;
  assign new_n12337_ = ~new_n5076_ & new_n12335_;
  assign new_n12338_ = ~new_n12336_ & ~new_n12337_;
  assign new_n12339_ = new_n4475_ & ~new_n12338_;
  assign new_n12340_ = lo0104 & new_n5083_;
  assign new_n12341_ = ~new_n12333_ & ~new_n12339_;
  assign new_n12342_ = ~new_n12340_ & new_n12341_;
  assign new_n12343_ = new_n3746_ & new_n12324_;
  assign new_n12344_ = ~new_n4096_ & new_n12325_;
  assign new_n12345_ = lo0104 & ~new_n12325_;
  assign new_n12346_ = ~new_n12344_ & ~new_n12345_;
  assign new_n12347_ = new_n5090_ & ~new_n12346_;
  assign new_n12348_ = ~new_n12343_ & ~new_n12347_;
  assign new_n12349_ = new_n5070_ & ~new_n12342_;
  assign new_n12350_ = new_n12348_ & ~new_n12349_;
  assign new_n12351_ = lo0104 & ~lo0841;
  assign new_n12352_ = new_n4020_ & new_n12325_;
  assign new_n12353_ = ~new_n5096_ & new_n12351_;
  assign new_n12354_ = ~new_n12352_ & ~new_n12353_;
  assign new_n12355_ = new_n12328_ & new_n12332_;
  assign new_n12356_ = new_n12350_ & new_n12355_;
  assign new_n12357_ = new_n12354_ & new_n12356_;
  assign new_n12358_ = new_n3804_ & new_n12325_;
  assign new_n12359_ = new_n3834_ & new_n12335_;
  assign new_n12360_ = new_n3678_ & new_n12359_;
  assign new_n12361_ = lo0104 & new_n5112_;
  assign new_n12362_ = new_n3810_ & new_n12351_;
  assign new_n12363_ = ~new_n12358_ & ~new_n12360_;
  assign new_n12364_ = ~new_n12361_ & new_n12363_;
  assign new_n12365_ = ~new_n12362_ & new_n12364_;
  assign new_n12366_ = ~new_n5105_ & new_n12351_;
  assign new_n12367_ = new_n12365_ & ~new_n12366_;
  assign new_n12368_ = new_n3815_ & new_n12324_;
  assign new_n12369_ = new_n4088_ & new_n12325_;
  assign new_n12370_ = ~new_n12368_ & ~new_n12369_;
  assign new_n12371_ = ~lo1044 & new_n12324_;
  assign new_n12372_ = new_n3820_ & new_n12351_;
  assign new_n12373_ = new_n3870_ & new_n12371_;
  assign new_n12374_ = ~new_n12372_ & ~new_n12373_;
  assign new_n12375_ = ~new_n4069_ & new_n12325_;
  assign new_n12376_ = new_n12367_ & new_n12370_;
  assign new_n12377_ = new_n12374_ & new_n12376_;
  assign new_n12378_ = ~new_n12375_ & new_n12377_;
  assign new_n12379_ = lo0104 & new_n5155_;
  assign new_n12380_ = new_n3777_ & new_n12379_;
  assign new_n12381_ = lo0104 & ~new_n4632_;
  assign new_n12382_ = new_n5565_ & new_n12381_;
  assign new_n12383_ = ~new_n12380_ & ~new_n12382_;
  assign new_n12384_ = ~new_n5460_ & new_n12324_;
  assign new_n12385_ = new_n12383_ & ~new_n12384_;
  assign new_n12386_ = lo0104 & new_n5562_;
  assign new_n12387_ = new_n4050_ & new_n12325_;
  assign new_n12388_ = new_n3763_ & new_n12351_;
  assign new_n12389_ = new_n3780_ & new_n12325_;
  assign new_n12390_ = ~new_n12388_ & ~new_n12389_;
  assign new_n12391_ = new_n3794_ & new_n12324_;
  assign new_n12392_ = new_n12390_ & ~new_n12391_;
  assign new_n12393_ = new_n12385_ & ~new_n12386_;
  assign new_n12394_ = ~new_n12387_ & new_n12393_;
  assign new_n12395_ = new_n12392_ & new_n12394_;
  assign new_n12396_ = new_n4041_ & new_n12325_;
  assign new_n12397_ = new_n12395_ & ~new_n12396_;
  assign new_n12398_ = lo0104 & new_n3678_;
  assign new_n12399_ = new_n3786_ & new_n12325_;
  assign new_n12400_ = new_n5139_ & new_n12398_;
  assign new_n12401_ = ~new_n12399_ & ~new_n12400_;
  assign new_n12402_ = new_n4007_ & new_n12371_;
  assign new_n12403_ = new_n3969_ & new_n12351_;
  assign new_n12404_ = ~new_n12402_ & ~new_n12403_;
  assign new_n12405_ = lo0104 & ~new_n5216_;
  assign new_n12406_ = new_n4133_ & new_n12325_;
  assign new_n12407_ = ~new_n12405_ & ~new_n12406_;
  assign new_n12408_ = new_n3974_ & new_n12335_;
  assign new_n12409_ = ~new_n4135_ & new_n12408_;
  assign new_n12410_ = lo0104 & new_n5225_;
  assign new_n12411_ = new_n12407_ & ~new_n12409_;
  assign new_n12412_ = ~new_n12410_ & new_n12411_;
  assign new_n12413_ = new_n3948_ & new_n12325_;
  assign new_n12414_ = new_n12412_ & ~new_n12413_;
  assign new_n12415_ = new_n12397_ & new_n12401_;
  assign new_n12416_ = new_n12404_ & new_n12415_;
  assign new_n12417_ = new_n12414_ & new_n12416_;
  assign new_n12418_ = lo0104 & new_n5194_;
  assign new_n12419_ = ~new_n12325_ & ~new_n12418_;
  assign new_n12420_ = new_n3936_ & ~new_n12419_;
  assign new_n12421_ = new_n3625_ & new_n12325_;
  assign new_n12422_ = ~new_n12420_ & ~new_n12421_;
  assign new_n12423_ = lo0104 & new_n3706_;
  assign new_n12424_ = lo0104 & new_n5608_;
  assign new_n12425_ = ~new_n5184_ & new_n12424_;
  assign new_n12426_ = new_n12422_ & ~new_n12423_;
  assign new_n12427_ = ~new_n12425_ & new_n12426_;
  assign new_n12428_ = ~new_n5201_ & new_n12351_;
  assign new_n12429_ = new_n12427_ & ~new_n12428_;
  assign new_n12430_ = ~lo0104 & new_n5230_;
  assign new_n12431_ = new_n4001_ & ~new_n12430_;
  assign new_n12432_ = lo0104 & new_n5135_;
  assign new_n12433_ = new_n12429_ & ~new_n12431_;
  assign new_n12434_ = ~new_n12432_ & new_n12433_;
  assign new_n12435_ = new_n12357_ & new_n12378_;
  assign new_n12436_ = new_n12417_ & new_n12435_;
  assign li0104 = ~new_n12434_ | ~new_n12436_;
  assign new_n12438_ = lo0106 & ~lo0841;
  assign new_n12439_ = ~new_n5201_ & new_n12438_;
  assign new_n12440_ = ~lo0024 & lo0106;
  assign new_n12441_ = lo0106 & new_n5194_;
  assign new_n12442_ = ~new_n12440_ & ~new_n12441_;
  assign new_n12443_ = new_n3936_ & ~new_n12442_;
  assign new_n12444_ = new_n3625_ & new_n12440_;
  assign new_n12445_ = ~new_n12443_ & ~new_n12444_;
  assign new_n12446_ = lo0106 & new_n5608_;
  assign new_n12447_ = ~new_n5184_ & new_n12446_;
  assign new_n12448_ = lo0106 & new_n3706_;
  assign new_n12449_ = ~new_n12439_ & new_n12445_;
  assign new_n12450_ = ~new_n12447_ & new_n12449_;
  assign new_n12451_ = ~new_n12448_ & new_n12450_;
  assign new_n12452_ = lo0106 & new_n5505_;
  assign new_n12453_ = lo0106 & ~new_n5216_;
  assign new_n12454_ = new_n4133_ & new_n12440_;
  assign new_n12455_ = ~new_n12453_ & ~new_n12454_;
  assign new_n12456_ = lo0106 & li0583;
  assign new_n12457_ = new_n3974_ & new_n12456_;
  assign new_n12458_ = ~new_n4135_ & new_n12457_;
  assign new_n12459_ = lo0106 & new_n5225_;
  assign new_n12460_ = new_n12455_ & ~new_n12458_;
  assign new_n12461_ = ~new_n12459_ & new_n12460_;
  assign new_n12462_ = new_n3948_ & new_n12440_;
  assign new_n12463_ = new_n12461_ & ~new_n12462_;
  assign new_n12464_ = lo0106 & ~lo0314;
  assign new_n12465_ = ~lo1044 & new_n12464_;
  assign new_n12466_ = new_n4007_ & new_n12465_;
  assign new_n12467_ = new_n3969_ & new_n12438_;
  assign new_n12468_ = ~new_n12466_ & ~new_n12467_;
  assign new_n12469_ = ~new_n12452_ & new_n12463_;
  assign new_n12470_ = new_n12468_ & new_n12469_;
  assign new_n12471_ = new_n12451_ & new_n12470_;
  assign new_n12472_ = new_n3985_ & new_n12464_;
  assign new_n12473_ = new_n4041_ & new_n12440_;
  assign new_n12474_ = ~new_n12472_ & ~new_n12473_;
  assign new_n12475_ = lo0106 & new_n5562_;
  assign new_n12476_ = new_n4050_ & new_n12440_;
  assign new_n12477_ = ~new_n12475_ & ~new_n12476_;
  assign new_n12478_ = new_n3763_ & new_n12438_;
  assign new_n12479_ = new_n3780_ & new_n12440_;
  assign new_n12480_ = ~new_n12478_ & ~new_n12479_;
  assign new_n12481_ = new_n3794_ & new_n12464_;
  assign new_n12482_ = new_n12480_ & ~new_n12481_;
  assign new_n12483_ = ~new_n5460_ & new_n12464_;
  assign new_n12484_ = lo0106 & ~new_n4632_;
  assign new_n12485_ = new_n5565_ & new_n12484_;
  assign new_n12486_ = lo0106 & new_n6643_;
  assign new_n12487_ = new_n12482_ & ~new_n12483_;
  assign new_n12488_ = ~new_n12485_ & new_n12487_;
  assign new_n12489_ = ~new_n12486_ & new_n12488_;
  assign new_n12490_ = new_n12477_ & new_n12489_;
  assign new_n12491_ = lo0106 & new_n5140_;
  assign new_n12492_ = new_n3786_ & new_n12440_;
  assign new_n12493_ = new_n12474_ & new_n12490_;
  assign new_n12494_ = ~new_n12491_ & new_n12493_;
  assign new_n12495_ = ~new_n12492_ & new_n12494_;
  assign new_n12496_ = new_n3979_ & new_n12464_;
  assign new_n12497_ = new_n12495_ & ~new_n12496_;
  assign new_n12498_ = lo0106 & ~lo0993;
  assign new_n12499_ = new_n3927_ & new_n12498_;
  assign new_n12500_ = new_n3940_ & new_n12440_;
  assign new_n12501_ = ~new_n12499_ & ~new_n12500_;
  assign new_n12502_ = lo0106 & new_n5135_;
  assign new_n12503_ = ~lo0024 & ~lo0106;
  assign new_n12504_ = new_n3953_ & ~new_n12503_;
  assign new_n12505_ = new_n12497_ & new_n12501_;
  assign new_n12506_ = ~new_n12502_ & new_n12505_;
  assign new_n12507_ = ~new_n12504_ & new_n12506_;
  assign new_n12508_ = new_n12471_ & new_n12507_;
  assign new_n12509_ = new_n3834_ & new_n12456_;
  assign new_n12510_ = new_n3678_ & new_n12509_;
  assign new_n12511_ = new_n3804_ & new_n12440_;
  assign new_n12512_ = ~new_n12510_ & ~new_n12511_;
  assign new_n12513_ = new_n3810_ & new_n12438_;
  assign new_n12514_ = lo0106 & new_n5112_;
  assign new_n12515_ = ~new_n12513_ & ~new_n12514_;
  assign new_n12516_ = new_n12512_ & new_n12515_;
  assign new_n12517_ = new_n4020_ & new_n12440_;
  assign new_n12518_ = ~new_n5096_ & new_n12438_;
  assign new_n12519_ = ~new_n12517_ & ~new_n12518_;
  assign new_n12520_ = ~new_n4096_ & new_n12440_;
  assign new_n12521_ = lo0106 & ~new_n12440_;
  assign new_n12522_ = ~new_n12520_ & ~new_n12521_;
  assign new_n12523_ = new_n5090_ & ~new_n12522_;
  assign new_n12524_ = new_n3746_ & new_n12464_;
  assign new_n12525_ = ~new_n12523_ & ~new_n12524_;
  assign new_n12526_ = lo0106 & new_n5071_;
  assign new_n12527_ = lo0106 & new_n4219_;
  assign new_n12528_ = ~new_n5074_ & new_n12527_;
  assign new_n12529_ = ~new_n5076_ & new_n12456_;
  assign new_n12530_ = ~new_n12528_ & ~new_n12529_;
  assign new_n12531_ = new_n4475_ & ~new_n12530_;
  assign new_n12532_ = lo0106 & new_n5083_;
  assign new_n12533_ = ~new_n12526_ & ~new_n12531_;
  assign new_n12534_ = ~new_n12532_ & new_n12533_;
  assign new_n12535_ = new_n5070_ & ~new_n12534_;
  assign new_n12536_ = new_n12516_ & new_n12519_;
  assign new_n12537_ = new_n12525_ & new_n12536_;
  assign new_n12538_ = ~new_n12535_ & new_n12537_;
  assign new_n12539_ = ~new_n5105_ & new_n12438_;
  assign new_n12540_ = new_n12538_ & ~new_n12539_;
  assign new_n12541_ = new_n3815_ & new_n12464_;
  assign new_n12542_ = new_n4088_ & new_n12440_;
  assign new_n12543_ = ~new_n12541_ & ~new_n12542_;
  assign new_n12544_ = new_n3820_ & new_n12438_;
  assign new_n12545_ = new_n3870_ & new_n12465_;
  assign new_n12546_ = ~new_n12544_ & ~new_n12545_;
  assign new_n12547_ = ~new_n4069_ & new_n12440_;
  assign new_n12548_ = new_n12546_ & ~new_n12547_;
  assign new_n12549_ = new_n12508_ & new_n12540_;
  assign new_n12550_ = new_n12543_ & new_n12549_;
  assign li0106 = ~new_n12548_ | ~new_n12550_;
  assign new_n12552_ = lo0107 & ~lo0841;
  assign new_n12553_ = ~new_n5201_ & new_n12552_;
  assign new_n12554_ = ~lo0024 & lo0107;
  assign new_n12555_ = lo0107 & new_n5194_;
  assign new_n12556_ = ~new_n12554_ & ~new_n12555_;
  assign new_n12557_ = new_n3936_ & ~new_n12556_;
  assign new_n12558_ = new_n3625_ & new_n12554_;
  assign new_n12559_ = ~new_n12557_ & ~new_n12558_;
  assign new_n12560_ = lo0107 & new_n5608_;
  assign new_n12561_ = ~new_n5184_ & new_n12560_;
  assign new_n12562_ = lo0107 & new_n3706_;
  assign new_n12563_ = ~new_n12553_ & new_n12559_;
  assign new_n12564_ = ~new_n12561_ & new_n12563_;
  assign new_n12565_ = ~new_n12562_ & new_n12564_;
  assign new_n12566_ = lo0107 & ~lo0314;
  assign new_n12567_ = ~new_n3940_ & ~new_n3953_;
  assign new_n12568_ = new_n12554_ & ~new_n12567_;
  assign new_n12569_ = new_n3979_ & new_n12566_;
  assign new_n12570_ = ~new_n12568_ & ~new_n12569_;
  assign new_n12571_ = new_n4050_ & new_n12554_;
  assign new_n12572_ = lo0107 & new_n5562_;
  assign new_n12573_ = lo0107 & new_n5155_;
  assign new_n12574_ = new_n3777_ & new_n12573_;
  assign new_n12575_ = lo0107 & ~new_n4632_;
  assign new_n12576_ = new_n5565_ & new_n12575_;
  assign new_n12577_ = ~new_n12574_ & ~new_n12576_;
  assign new_n12578_ = ~new_n5460_ & new_n12566_;
  assign new_n12579_ = new_n12577_ & ~new_n12578_;
  assign new_n12580_ = new_n3763_ & new_n12552_;
  assign new_n12581_ = new_n3780_ & new_n12554_;
  assign new_n12582_ = ~new_n12580_ & ~new_n12581_;
  assign new_n12583_ = new_n3794_ & new_n12566_;
  assign new_n12584_ = new_n12582_ & ~new_n12583_;
  assign new_n12585_ = ~new_n12571_ & ~new_n12572_;
  assign new_n12586_ = new_n12579_ & new_n12585_;
  assign new_n12587_ = new_n12584_ & new_n12586_;
  assign new_n12588_ = lo0107 & new_n5140_;
  assign new_n12589_ = new_n3786_ & new_n12554_;
  assign new_n12590_ = ~new_n12588_ & ~new_n12589_;
  assign new_n12591_ = new_n12587_ & new_n12590_;
  assign new_n12592_ = new_n3985_ & new_n12566_;
  assign new_n12593_ = new_n4041_ & new_n12554_;
  assign new_n12594_ = ~new_n12592_ & ~new_n12593_;
  assign new_n12595_ = new_n12570_ & new_n12591_;
  assign new_n12596_ = new_n12594_ & new_n12595_;
  assign new_n12597_ = new_n12565_ & new_n12596_;
  assign new_n12598_ = lo0107 & new_n5505_;
  assign new_n12599_ = lo0107 & ~new_n5216_;
  assign new_n12600_ = new_n4133_ & new_n12554_;
  assign new_n12601_ = ~new_n12599_ & ~new_n12600_;
  assign new_n12602_ = lo0107 & li0583;
  assign new_n12603_ = new_n3974_ & new_n12602_;
  assign new_n12604_ = ~new_n4135_ & new_n12603_;
  assign new_n12605_ = lo0107 & new_n5225_;
  assign new_n12606_ = new_n12601_ & ~new_n12604_;
  assign new_n12607_ = ~new_n12605_ & new_n12606_;
  assign new_n12608_ = new_n3948_ & new_n12554_;
  assign new_n12609_ = new_n12607_ & ~new_n12608_;
  assign new_n12610_ = ~lo1044 & new_n12566_;
  assign new_n12611_ = new_n4007_ & new_n12610_;
  assign new_n12612_ = new_n3969_ & new_n12552_;
  assign new_n12613_ = ~new_n12611_ & ~new_n12612_;
  assign new_n12614_ = new_n12609_ & new_n12613_;
  assign new_n12615_ = lo0107 & new_n5135_;
  assign new_n12616_ = ~lo0107 & ~lo0993;
  assign new_n12617_ = new_n3927_ & ~new_n12616_;
  assign new_n12618_ = ~new_n12598_ & new_n12614_;
  assign new_n12619_ = ~new_n12615_ & new_n12618_;
  assign new_n12620_ = ~new_n12617_ & new_n12619_;
  assign new_n12621_ = new_n12597_ & new_n12620_;
  assign new_n12622_ = new_n3834_ & new_n12602_;
  assign new_n12623_ = new_n3678_ & new_n12622_;
  assign new_n12624_ = new_n3804_ & new_n12554_;
  assign new_n12625_ = ~new_n12623_ & ~new_n12624_;
  assign new_n12626_ = new_n3810_ & new_n12552_;
  assign new_n12627_ = lo0107 & new_n5112_;
  assign new_n12628_ = ~new_n12626_ & ~new_n12627_;
  assign new_n12629_ = new_n12625_ & new_n12628_;
  assign new_n12630_ = new_n4020_ & new_n12554_;
  assign new_n12631_ = ~new_n5096_ & new_n12552_;
  assign new_n12632_ = ~new_n12630_ & ~new_n12631_;
  assign new_n12633_ = ~new_n4096_ & new_n12554_;
  assign new_n12634_ = lo0107 & ~new_n12554_;
  assign new_n12635_ = ~new_n12633_ & ~new_n12634_;
  assign new_n12636_ = new_n5090_ & ~new_n12635_;
  assign new_n12637_ = new_n3746_ & new_n12566_;
  assign new_n12638_ = ~new_n12636_ & ~new_n12637_;
  assign new_n12639_ = lo0107 & new_n5071_;
  assign new_n12640_ = lo0107 & new_n4219_;
  assign new_n12641_ = ~new_n5074_ & new_n12640_;
  assign new_n12642_ = ~new_n5076_ & new_n12602_;
  assign new_n12643_ = ~new_n12641_ & ~new_n12642_;
  assign new_n12644_ = new_n4475_ & ~new_n12643_;
  assign new_n12645_ = lo0107 & new_n5083_;
  assign new_n12646_ = ~new_n12639_ & ~new_n12644_;
  assign new_n12647_ = ~new_n12645_ & new_n12646_;
  assign new_n12648_ = new_n5070_ & ~new_n12647_;
  assign new_n12649_ = new_n12629_ & new_n12632_;
  assign new_n12650_ = new_n12638_ & new_n12649_;
  assign new_n12651_ = ~new_n12648_ & new_n12650_;
  assign new_n12652_ = ~new_n5105_ & new_n12552_;
  assign new_n12653_ = new_n12651_ & ~new_n12652_;
  assign new_n12654_ = new_n3815_ & new_n12566_;
  assign new_n12655_ = new_n4088_ & new_n12554_;
  assign new_n12656_ = ~new_n12654_ & ~new_n12655_;
  assign new_n12657_ = new_n3820_ & new_n12552_;
  assign new_n12658_ = new_n3870_ & new_n12610_;
  assign new_n12659_ = ~new_n12657_ & ~new_n12658_;
  assign new_n12660_ = ~new_n4069_ & new_n12554_;
  assign new_n12661_ = new_n12659_ & ~new_n12660_;
  assign new_n12662_ = new_n12621_ & new_n12653_;
  assign new_n12663_ = new_n12656_ & new_n12662_;
  assign li0107 = ~new_n12661_ | ~new_n12663_;
  assign new_n12665_ = lo0108 & ~lo0841;
  assign new_n12666_ = ~lo0024 & lo0108;
  assign new_n12667_ = new_n3804_ & new_n12666_;
  assign new_n12668_ = lo0108 & li0583;
  assign new_n12669_ = new_n3834_ & new_n12668_;
  assign new_n12670_ = new_n3678_ & new_n12669_;
  assign new_n12671_ = lo0108 & new_n5112_;
  assign new_n12672_ = new_n3810_ & new_n12665_;
  assign new_n12673_ = ~new_n12667_ & ~new_n12670_;
  assign new_n12674_ = ~new_n12671_ & new_n12673_;
  assign new_n12675_ = ~new_n12672_ & new_n12674_;
  assign new_n12676_ = ~new_n5105_ & new_n12665_;
  assign new_n12677_ = new_n12675_ & ~new_n12676_;
  assign new_n12678_ = lo0108 & ~lo0314;
  assign new_n12679_ = new_n3815_ & new_n12678_;
  assign new_n12680_ = new_n4088_ & new_n12666_;
  assign new_n12681_ = ~new_n12679_ & ~new_n12680_;
  assign new_n12682_ = ~lo1044 & new_n12678_;
  assign new_n12683_ = new_n3820_ & new_n12665_;
  assign new_n12684_ = new_n3870_ & new_n12682_;
  assign new_n12685_ = ~new_n12683_ & ~new_n12684_;
  assign new_n12686_ = ~new_n4069_ & new_n12666_;
  assign new_n12687_ = new_n12677_ & new_n12681_;
  assign new_n12688_ = new_n12685_ & new_n12687_;
  assign new_n12689_ = ~new_n12686_ & new_n12688_;
  assign new_n12690_ = new_n3763_ & new_n12665_;
  assign new_n12691_ = new_n3780_ & new_n12666_;
  assign new_n12692_ = ~new_n12690_ & ~new_n12691_;
  assign new_n12693_ = new_n3794_ & new_n12678_;
  assign new_n12694_ = new_n12692_ & ~new_n12693_;
  assign new_n12695_ = ~new_n5460_ & new_n12678_;
  assign new_n12696_ = lo0108 & ~new_n4632_;
  assign new_n12697_ = new_n5565_ & new_n12696_;
  assign new_n12698_ = lo0108 & new_n6643_;
  assign new_n12699_ = new_n12694_ & ~new_n12695_;
  assign new_n12700_ = ~new_n12697_ & new_n12699_;
  assign new_n12701_ = ~new_n12698_ & new_n12700_;
  assign new_n12702_ = lo0108 & new_n5671_;
  assign new_n12703_ = new_n3940_ & new_n12666_;
  assign new_n12704_ = ~new_n12702_ & ~new_n12703_;
  assign new_n12705_ = new_n12701_ & new_n12704_;
  assign new_n12706_ = new_n12689_ & new_n12705_;
  assign new_n12707_ = lo0108 & new_n5071_;
  assign new_n12708_ = lo0108 & new_n4219_;
  assign new_n12709_ = ~new_n5074_ & new_n12708_;
  assign new_n12710_ = ~new_n5076_ & new_n12668_;
  assign new_n12711_ = ~new_n12709_ & ~new_n12710_;
  assign new_n12712_ = new_n4475_ & ~new_n12711_;
  assign new_n12713_ = lo0108 & new_n5083_;
  assign new_n12714_ = ~new_n12707_ & ~new_n12712_;
  assign new_n12715_ = ~new_n12713_ & new_n12714_;
  assign new_n12716_ = new_n3746_ & new_n12678_;
  assign new_n12717_ = ~new_n4096_ & new_n12666_;
  assign new_n12718_ = lo0108 & ~new_n12666_;
  assign new_n12719_ = ~new_n12717_ & ~new_n12718_;
  assign new_n12720_ = new_n5090_ & ~new_n12719_;
  assign new_n12721_ = ~new_n12716_ & ~new_n12720_;
  assign new_n12722_ = new_n5070_ & ~new_n12715_;
  assign new_n12723_ = new_n12721_ & ~new_n12722_;
  assign new_n12724_ = new_n4007_ & new_n12682_;
  assign new_n12725_ = new_n3969_ & new_n12665_;
  assign new_n12726_ = ~new_n12724_ & ~new_n12725_;
  assign new_n12727_ = new_n3948_ & new_n12666_;
  assign new_n12728_ = new_n3974_ & new_n12668_;
  assign new_n12729_ = ~new_n4135_ & new_n12728_;
  assign new_n12730_ = lo0108 & new_n5225_;
  assign new_n12731_ = ~new_n12729_ & ~new_n12730_;
  assign new_n12732_ = lo0108 & ~new_n5216_;
  assign new_n12733_ = new_n4133_ & new_n12666_;
  assign new_n12734_ = ~new_n12732_ & ~new_n12733_;
  assign new_n12735_ = new_n12726_ & ~new_n12727_;
  assign new_n12736_ = new_n12731_ & new_n12735_;
  assign new_n12737_ = new_n12734_ & new_n12736_;
  assign new_n12738_ = new_n3985_ & new_n12678_;
  assign new_n12739_ = new_n12737_ & ~new_n12738_;
  assign new_n12740_ = new_n12723_ & new_n12739_;
  assign new_n12741_ = new_n4020_ & new_n12666_;
  assign new_n12742_ = ~new_n5096_ & new_n12665_;
  assign new_n12743_ = ~new_n12741_ & ~new_n12742_;
  assign new_n12744_ = new_n3979_ & new_n12678_;
  assign new_n12745_ = new_n3953_ & new_n12666_;
  assign new_n12746_ = ~new_n12744_ & ~new_n12745_;
  assign new_n12747_ = new_n12743_ & new_n12746_;
  assign new_n12748_ = ~new_n3959_ & new_n12747_;
  assign new_n12749_ = ~new_n3989_ & new_n12748_;
  assign new_n12750_ = lo0108 & new_n5505_;
  assign new_n12751_ = new_n12749_ & ~new_n12750_;
  assign new_n12752_ = new_n12740_ & new_n12751_;
  assign new_n12753_ = lo0108 & new_n5562_;
  assign new_n12754_ = new_n4050_ & new_n12666_;
  assign new_n12755_ = ~new_n12753_ & ~new_n12754_;
  assign new_n12756_ = new_n4041_ & new_n12666_;
  assign new_n12757_ = new_n12755_ & ~new_n12756_;
  assign new_n12758_ = lo0108 & new_n5140_;
  assign new_n12759_ = new_n3786_ & new_n12666_;
  assign new_n12760_ = ~new_n3769_ & new_n12757_;
  assign new_n12761_ = ~new_n12758_ & new_n12760_;
  assign new_n12762_ = ~new_n12759_ & new_n12761_;
  assign new_n12763_ = lo0108 & ~new_n5134_;
  assign new_n12764_ = new_n5133_ & new_n12763_;
  assign new_n12765_ = new_n12762_ & ~new_n12764_;
  assign new_n12766_ = ~new_n5201_ & new_n12665_;
  assign new_n12767_ = lo0108 & new_n5194_;
  assign new_n12768_ = ~new_n12666_ & ~new_n12767_;
  assign new_n12769_ = new_n3936_ & ~new_n12768_;
  assign new_n12770_ = new_n3625_ & new_n12666_;
  assign new_n12771_ = ~new_n12769_ & ~new_n12770_;
  assign new_n12772_ = lo0108 & new_n5608_;
  assign new_n12773_ = ~new_n5184_ & new_n12772_;
  assign new_n12774_ = lo0108 & new_n3706_;
  assign new_n12775_ = ~new_n12766_ & new_n12771_;
  assign new_n12776_ = ~new_n12773_ & new_n12775_;
  assign new_n12777_ = ~new_n12774_ & new_n12776_;
  assign new_n12778_ = new_n12706_ & new_n12752_;
  assign new_n12779_ = new_n12765_ & new_n12778_;
  assign li0108 = ~new_n12777_ | ~new_n12779_;
  assign new_n12781_ = lo0109 & ~lo0841;
  assign new_n12782_ = ~new_n5201_ & new_n12781_;
  assign new_n12783_ = ~lo0024 & lo0109;
  assign new_n12784_ = lo0109 & new_n5194_;
  assign new_n12785_ = ~new_n12783_ & ~new_n12784_;
  assign new_n12786_ = new_n3936_ & ~new_n12785_;
  assign new_n12787_ = new_n3625_ & new_n12783_;
  assign new_n12788_ = ~new_n12786_ & ~new_n12787_;
  assign new_n12789_ = lo0109 & new_n5608_;
  assign new_n12790_ = ~new_n5184_ & new_n12789_;
  assign new_n12791_ = lo0109 & new_n3706_;
  assign new_n12792_ = ~new_n12782_ & new_n12788_;
  assign new_n12793_ = ~new_n12790_ & new_n12792_;
  assign new_n12794_ = ~new_n12791_ & new_n12793_;
  assign new_n12795_ = lo0109 & new_n5505_;
  assign new_n12796_ = lo0109 & ~new_n5216_;
  assign new_n12797_ = new_n4133_ & new_n12783_;
  assign new_n12798_ = ~new_n12796_ & ~new_n12797_;
  assign new_n12799_ = lo0109 & li0583;
  assign new_n12800_ = new_n3974_ & new_n12799_;
  assign new_n12801_ = ~new_n4135_ & new_n12800_;
  assign new_n12802_ = lo0109 & new_n5225_;
  assign new_n12803_ = new_n12798_ & ~new_n12801_;
  assign new_n12804_ = ~new_n12802_ & new_n12803_;
  assign new_n12805_ = new_n3948_ & new_n12783_;
  assign new_n12806_ = new_n12804_ & ~new_n12805_;
  assign new_n12807_ = lo0109 & ~lo0314;
  assign new_n12808_ = ~lo1044 & new_n12807_;
  assign new_n12809_ = new_n4007_ & new_n12808_;
  assign new_n12810_ = new_n3969_ & new_n12781_;
  assign new_n12811_ = ~new_n12809_ & ~new_n12810_;
  assign new_n12812_ = ~new_n12795_ & new_n12806_;
  assign new_n12813_ = new_n12811_ & new_n12812_;
  assign new_n12814_ = new_n12794_ & new_n12813_;
  assign new_n12815_ = new_n3985_ & new_n12807_;
  assign new_n12816_ = new_n4041_ & new_n12783_;
  assign new_n12817_ = ~new_n12815_ & ~new_n12816_;
  assign new_n12818_ = lo0109 & new_n5562_;
  assign new_n12819_ = new_n4050_ & new_n12783_;
  assign new_n12820_ = ~new_n12818_ & ~new_n12819_;
  assign new_n12821_ = new_n3763_ & new_n12781_;
  assign new_n12822_ = new_n3780_ & new_n12783_;
  assign new_n12823_ = ~new_n12821_ & ~new_n12822_;
  assign new_n12824_ = new_n3794_ & new_n12807_;
  assign new_n12825_ = new_n12823_ & ~new_n12824_;
  assign new_n12826_ = ~new_n5460_ & new_n12807_;
  assign new_n12827_ = lo0109 & ~new_n4632_;
  assign new_n12828_ = new_n5565_ & new_n12827_;
  assign new_n12829_ = lo0109 & new_n6643_;
  assign new_n12830_ = new_n12825_ & ~new_n12826_;
  assign new_n12831_ = ~new_n12828_ & new_n12830_;
  assign new_n12832_ = ~new_n12829_ & new_n12831_;
  assign new_n12833_ = new_n12820_ & new_n12832_;
  assign new_n12834_ = lo0109 & new_n5140_;
  assign new_n12835_ = new_n3786_ & new_n12783_;
  assign new_n12836_ = new_n12817_ & new_n12833_;
  assign new_n12837_ = ~new_n12834_ & new_n12836_;
  assign new_n12838_ = ~new_n12835_ & new_n12837_;
  assign new_n12839_ = new_n3940_ & new_n12783_;
  assign new_n12840_ = new_n12838_ & ~new_n12839_;
  assign new_n12841_ = lo0109 & ~lo0993;
  assign new_n12842_ = new_n3927_ & new_n12841_;
  assign new_n12843_ = new_n3953_ & new_n12783_;
  assign new_n12844_ = ~new_n12842_ & ~new_n12843_;
  assign new_n12845_ = lo0314 & new_n3979_;
  assign new_n12846_ = lo0109 & ~new_n5134_;
  assign new_n12847_ = new_n5133_ & new_n12846_;
  assign new_n12848_ = lo0109 & new_n3979_;
  assign new_n12849_ = ~new_n12847_ & ~new_n12848_;
  assign new_n12850_ = new_n12840_ & new_n12844_;
  assign new_n12851_ = ~new_n12845_ & new_n12850_;
  assign new_n12852_ = new_n12849_ & new_n12851_;
  assign new_n12853_ = new_n12814_ & new_n12852_;
  assign new_n12854_ = new_n3834_ & new_n12799_;
  assign new_n12855_ = new_n3678_ & new_n12854_;
  assign new_n12856_ = new_n3804_ & new_n12783_;
  assign new_n12857_ = ~new_n12855_ & ~new_n12856_;
  assign new_n12858_ = new_n3810_ & new_n12781_;
  assign new_n12859_ = lo0109 & new_n5112_;
  assign new_n12860_ = ~new_n12858_ & ~new_n12859_;
  assign new_n12861_ = new_n12857_ & new_n12860_;
  assign new_n12862_ = new_n4020_ & new_n12783_;
  assign new_n12863_ = ~new_n5096_ & new_n12781_;
  assign new_n12864_ = ~new_n12862_ & ~new_n12863_;
  assign new_n12865_ = ~new_n4096_ & new_n12783_;
  assign new_n12866_ = lo0109 & ~new_n12783_;
  assign new_n12867_ = ~new_n12865_ & ~new_n12866_;
  assign new_n12868_ = new_n5090_ & ~new_n12867_;
  assign new_n12869_ = new_n3746_ & new_n12807_;
  assign new_n12870_ = ~new_n12868_ & ~new_n12869_;
  assign new_n12871_ = lo0109 & new_n5071_;
  assign new_n12872_ = lo0109 & new_n4219_;
  assign new_n12873_ = ~new_n5074_ & new_n12872_;
  assign new_n12874_ = ~new_n5076_ & new_n12799_;
  assign new_n12875_ = ~new_n12873_ & ~new_n12874_;
  assign new_n12876_ = new_n4475_ & ~new_n12875_;
  assign new_n12877_ = lo0109 & new_n5083_;
  assign new_n12878_ = ~new_n12871_ & ~new_n12876_;
  assign new_n12879_ = ~new_n12877_ & new_n12878_;
  assign new_n12880_ = new_n5070_ & ~new_n12879_;
  assign new_n12881_ = new_n12861_ & new_n12864_;
  assign new_n12882_ = new_n12870_ & new_n12881_;
  assign new_n12883_ = ~new_n12880_ & new_n12882_;
  assign new_n12884_ = ~new_n5105_ & new_n12781_;
  assign new_n12885_ = new_n12883_ & ~new_n12884_;
  assign new_n12886_ = new_n3815_ & new_n12807_;
  assign new_n12887_ = new_n4088_ & new_n12783_;
  assign new_n12888_ = ~new_n12886_ & ~new_n12887_;
  assign new_n12889_ = new_n3820_ & new_n12781_;
  assign new_n12890_ = new_n3870_ & new_n12808_;
  assign new_n12891_ = ~new_n12889_ & ~new_n12890_;
  assign new_n12892_ = ~new_n4069_ & new_n12783_;
  assign new_n12893_ = new_n12891_ & ~new_n12892_;
  assign new_n12894_ = new_n12853_ & new_n12885_;
  assign new_n12895_ = new_n12888_ & new_n12894_;
  assign li0109 = ~new_n12893_ | ~new_n12895_;
  assign new_n12897_ = lo0110 & ~lo0841;
  assign new_n12898_ = ~new_n5201_ & new_n12897_;
  assign new_n12899_ = ~lo0024 & lo0110;
  assign new_n12900_ = lo0110 & new_n5194_;
  assign new_n12901_ = ~new_n12899_ & ~new_n12900_;
  assign new_n12902_ = new_n3936_ & ~new_n12901_;
  assign new_n12903_ = new_n3625_ & new_n12899_;
  assign new_n12904_ = ~new_n12902_ & ~new_n12903_;
  assign new_n12905_ = lo0110 & new_n7163_;
  assign new_n12906_ = lo0110 & new_n3706_;
  assign new_n12907_ = ~new_n12898_ & new_n12904_;
  assign new_n12908_ = ~new_n12905_ & new_n12907_;
  assign new_n12909_ = ~new_n12906_ & new_n12908_;
  assign new_n12910_ = lo0110 & new_n5505_;
  assign new_n12911_ = lo0110 & ~new_n5216_;
  assign new_n12912_ = new_n4133_ & new_n12899_;
  assign new_n12913_ = ~new_n12911_ & ~new_n12912_;
  assign new_n12914_ = lo0110 & li0583;
  assign new_n12915_ = new_n3974_ & new_n12914_;
  assign new_n12916_ = ~new_n4135_ & new_n12915_;
  assign new_n12917_ = lo0110 & new_n5225_;
  assign new_n12918_ = new_n12913_ & ~new_n12916_;
  assign new_n12919_ = ~new_n12917_ & new_n12918_;
  assign new_n12920_ = new_n3948_ & new_n12899_;
  assign new_n12921_ = new_n12919_ & ~new_n12920_;
  assign new_n12922_ = lo0110 & ~lo0314;
  assign new_n12923_ = ~lo1044 & new_n12922_;
  assign new_n12924_ = new_n4007_ & new_n12923_;
  assign new_n12925_ = new_n3969_ & new_n12897_;
  assign new_n12926_ = ~new_n12924_ & ~new_n12925_;
  assign new_n12927_ = ~new_n12910_ & new_n12921_;
  assign new_n12928_ = new_n12926_ & new_n12927_;
  assign new_n12929_ = new_n12909_ & new_n12928_;
  assign new_n12930_ = new_n3979_ & new_n12922_;
  assign new_n12931_ = new_n4041_ & new_n12899_;
  assign new_n12932_ = ~new_n12930_ & ~new_n12931_;
  assign new_n12933_ = lo0110 & new_n5562_;
  assign new_n12934_ = new_n4050_ & new_n12899_;
  assign new_n12935_ = ~new_n12933_ & ~new_n12934_;
  assign new_n12936_ = new_n3763_ & new_n12897_;
  assign new_n12937_ = new_n3780_ & new_n12899_;
  assign new_n12938_ = ~new_n12936_ & ~new_n12937_;
  assign new_n12939_ = new_n3794_ & new_n12922_;
  assign new_n12940_ = new_n12938_ & ~new_n12939_;
  assign new_n12941_ = ~new_n5460_ & new_n12922_;
  assign new_n12942_ = lo0110 & ~new_n4632_;
  assign new_n12943_ = new_n5565_ & new_n12942_;
  assign new_n12944_ = lo0110 & new_n6643_;
  assign new_n12945_ = new_n12940_ & ~new_n12941_;
  assign new_n12946_ = ~new_n12943_ & new_n12945_;
  assign new_n12947_ = ~new_n12944_ & new_n12946_;
  assign new_n12948_ = new_n12935_ & new_n12947_;
  assign new_n12949_ = lo0110 & new_n5140_;
  assign new_n12950_ = new_n3786_ & new_n12899_;
  assign new_n12951_ = new_n12932_ & new_n12948_;
  assign new_n12952_ = ~new_n12949_ & new_n12951_;
  assign new_n12953_ = ~new_n12950_ & new_n12952_;
  assign new_n12954_ = new_n3940_ & new_n12899_;
  assign new_n12955_ = new_n12953_ & ~new_n12954_;
  assign new_n12956_ = lo0110 & ~lo0993;
  assign new_n12957_ = new_n3927_ & new_n12956_;
  assign new_n12958_ = new_n3953_ & new_n12899_;
  assign new_n12959_ = ~new_n12957_ & ~new_n12958_;
  assign new_n12960_ = lo0110 & new_n5135_;
  assign new_n12961_ = ~lo0110 & ~lo0314;
  assign new_n12962_ = new_n3985_ & ~new_n12961_;
  assign new_n12963_ = new_n12955_ & new_n12959_;
  assign new_n12964_ = ~new_n12960_ & new_n12963_;
  assign new_n12965_ = ~new_n12962_ & new_n12964_;
  assign new_n12966_ = new_n12929_ & new_n12965_;
  assign new_n12967_ = new_n3834_ & new_n12914_;
  assign new_n12968_ = new_n3678_ & new_n12967_;
  assign new_n12969_ = new_n3804_ & new_n12899_;
  assign new_n12970_ = ~new_n12968_ & ~new_n12969_;
  assign new_n12971_ = new_n3810_ & new_n12897_;
  assign new_n12972_ = lo0110 & new_n5112_;
  assign new_n12973_ = ~new_n12971_ & ~new_n12972_;
  assign new_n12974_ = new_n12970_ & new_n12973_;
  assign new_n12975_ = new_n4020_ & new_n12899_;
  assign new_n12976_ = ~new_n5096_ & new_n12897_;
  assign new_n12977_ = ~new_n12975_ & ~new_n12976_;
  assign new_n12978_ = ~new_n4096_ & new_n12899_;
  assign new_n12979_ = lo0110 & ~new_n12899_;
  assign new_n12980_ = ~new_n12978_ & ~new_n12979_;
  assign new_n12981_ = new_n5090_ & ~new_n12980_;
  assign new_n12982_ = new_n3746_ & new_n12922_;
  assign new_n12983_ = ~new_n12981_ & ~new_n12982_;
  assign new_n12984_ = lo0110 & new_n5071_;
  assign new_n12985_ = lo0110 & new_n4219_;
  assign new_n12986_ = ~new_n5074_ & new_n12985_;
  assign new_n12987_ = ~new_n5076_ & new_n12914_;
  assign new_n12988_ = ~new_n12986_ & ~new_n12987_;
  assign new_n12989_ = new_n4475_ & ~new_n12988_;
  assign new_n12990_ = lo0110 & new_n5083_;
  assign new_n12991_ = ~new_n12984_ & ~new_n12989_;
  assign new_n12992_ = ~new_n12990_ & new_n12991_;
  assign new_n12993_ = new_n5070_ & ~new_n12992_;
  assign new_n12994_ = new_n12974_ & new_n12977_;
  assign new_n12995_ = new_n12983_ & new_n12994_;
  assign new_n12996_ = ~new_n12993_ & new_n12995_;
  assign new_n12997_ = ~new_n5105_ & new_n12897_;
  assign new_n12998_ = new_n12996_ & ~new_n12997_;
  assign new_n12999_ = new_n3815_ & new_n12922_;
  assign new_n13000_ = new_n4088_ & new_n12899_;
  assign new_n13001_ = ~new_n12999_ & ~new_n13000_;
  assign new_n13002_ = new_n3820_ & new_n12897_;
  assign new_n13003_ = new_n3870_ & new_n12923_;
  assign new_n13004_ = ~new_n13002_ & ~new_n13003_;
  assign new_n13005_ = ~new_n4069_ & new_n12899_;
  assign new_n13006_ = new_n13004_ & ~new_n13005_;
  assign new_n13007_ = new_n12966_ & new_n12998_;
  assign new_n13008_ = new_n13001_ & new_n13007_;
  assign li0110 = ~new_n13006_ | ~new_n13008_;
  assign new_n13010_ = lo0111 & ~lo0841;
  assign new_n13011_ = ~new_n5201_ & new_n13010_;
  assign new_n13012_ = ~lo0024 & lo0111;
  assign new_n13013_ = lo0111 & new_n5194_;
  assign new_n13014_ = ~new_n13012_ & ~new_n13013_;
  assign new_n13015_ = new_n3936_ & ~new_n13014_;
  assign new_n13016_ = new_n3625_ & new_n13012_;
  assign new_n13017_ = ~new_n13015_ & ~new_n13016_;
  assign new_n13018_ = lo0111 & new_n5818_;
  assign new_n13019_ = ~new_n5184_ & new_n13018_;
  assign new_n13020_ = lo0111 & new_n3706_;
  assign new_n13021_ = ~new_n13011_ & new_n13017_;
  assign new_n13022_ = ~new_n13019_ & new_n13021_;
  assign new_n13023_ = ~new_n13020_ & new_n13022_;
  assign new_n13024_ = lo0111 & new_n5505_;
  assign new_n13025_ = lo0111 & ~new_n5216_;
  assign new_n13026_ = new_n4133_ & new_n13012_;
  assign new_n13027_ = ~new_n13025_ & ~new_n13026_;
  assign new_n13028_ = lo0111 & li0583;
  assign new_n13029_ = new_n3974_ & new_n13028_;
  assign new_n13030_ = ~new_n4135_ & new_n13029_;
  assign new_n13031_ = lo0111 & new_n5225_;
  assign new_n13032_ = new_n13027_ & ~new_n13030_;
  assign new_n13033_ = ~new_n13031_ & new_n13032_;
  assign new_n13034_ = new_n3948_ & new_n13012_;
  assign new_n13035_ = new_n13033_ & ~new_n13034_;
  assign new_n13036_ = lo0111 & ~lo0314;
  assign new_n13037_ = ~lo1044 & new_n13036_;
  assign new_n13038_ = new_n4007_ & new_n13037_;
  assign new_n13039_ = new_n3969_ & new_n13010_;
  assign new_n13040_ = ~new_n13038_ & ~new_n13039_;
  assign new_n13041_ = ~new_n13024_ & new_n13035_;
  assign new_n13042_ = new_n13040_ & new_n13041_;
  assign new_n13043_ = new_n13023_ & new_n13042_;
  assign new_n13044_ = lo0111 & new_n5562_;
  assign new_n13045_ = new_n4050_ & new_n13012_;
  assign new_n13046_ = ~new_n13044_ & ~new_n13045_;
  assign new_n13047_ = new_n3763_ & new_n13010_;
  assign new_n13048_ = new_n3780_ & new_n13012_;
  assign new_n13049_ = ~new_n13047_ & ~new_n13048_;
  assign new_n13050_ = new_n3794_ & new_n13036_;
  assign new_n13051_ = new_n13049_ & ~new_n13050_;
  assign new_n13052_ = ~new_n5460_ & new_n13036_;
  assign new_n13053_ = lo0111 & ~new_n4632_;
  assign new_n13054_ = new_n5565_ & new_n13053_;
  assign new_n13055_ = lo0111 & new_n6643_;
  assign new_n13056_ = new_n13051_ & ~new_n13052_;
  assign new_n13057_ = ~new_n13054_ & new_n13056_;
  assign new_n13058_ = ~new_n13055_ & new_n13057_;
  assign new_n13059_ = new_n13046_ & new_n13058_;
  assign new_n13060_ = new_n3786_ & new_n13012_;
  assign new_n13061_ = lo0111 & new_n5140_;
  assign new_n13062_ = new_n3953_ & new_n13012_;
  assign new_n13063_ = new_n3979_ & new_n13036_;
  assign new_n13064_ = ~new_n13062_ & ~new_n13063_;
  assign new_n13065_ = ~new_n13060_ & ~new_n13061_;
  assign new_n13066_ = new_n13064_ & new_n13065_;
  assign new_n13067_ = lo0111 & new_n5133_;
  assign new_n13068_ = ~new_n5134_ & new_n13067_;
  assign new_n13069_ = lo0111 & ~lo0993;
  assign new_n13070_ = ~lo0024 & ~lo0111;
  assign new_n13071_ = new_n3927_ & new_n13069_;
  assign new_n13072_ = new_n3940_ & ~new_n13070_;
  assign new_n13073_ = ~new_n13071_ & ~new_n13072_;
  assign new_n13074_ = ~new_n13068_ & new_n13073_;
  assign new_n13075_ = new_n13066_ & new_n13074_;
  assign new_n13076_ = new_n3985_ & new_n13036_;
  assign new_n13077_ = new_n4041_ & new_n13012_;
  assign new_n13078_ = ~new_n13076_ & ~new_n13077_;
  assign new_n13079_ = new_n13059_ & new_n13075_;
  assign new_n13080_ = new_n13078_ & new_n13079_;
  assign new_n13081_ = new_n13043_ & new_n13080_;
  assign new_n13082_ = new_n3834_ & new_n13028_;
  assign new_n13083_ = new_n3678_ & new_n13082_;
  assign new_n13084_ = new_n3804_ & new_n13012_;
  assign new_n13085_ = ~new_n13083_ & ~new_n13084_;
  assign new_n13086_ = new_n3810_ & new_n13010_;
  assign new_n13087_ = lo0111 & new_n5112_;
  assign new_n13088_ = ~new_n13086_ & ~new_n13087_;
  assign new_n13089_ = new_n13085_ & new_n13088_;
  assign new_n13090_ = new_n4020_ & new_n13012_;
  assign new_n13091_ = ~new_n5096_ & new_n13010_;
  assign new_n13092_ = ~new_n13090_ & ~new_n13091_;
  assign new_n13093_ = ~new_n4096_ & new_n13012_;
  assign new_n13094_ = lo0111 & ~new_n13012_;
  assign new_n13095_ = ~new_n13093_ & ~new_n13094_;
  assign new_n13096_ = new_n5090_ & ~new_n13095_;
  assign new_n13097_ = new_n3746_ & new_n13036_;
  assign new_n13098_ = ~new_n13096_ & ~new_n13097_;
  assign new_n13099_ = lo0111 & new_n5071_;
  assign new_n13100_ = lo0111 & new_n4219_;
  assign new_n13101_ = ~new_n5074_ & new_n13100_;
  assign new_n13102_ = ~new_n5076_ & new_n13028_;
  assign new_n13103_ = ~new_n13101_ & ~new_n13102_;
  assign new_n13104_ = new_n4475_ & ~new_n13103_;
  assign new_n13105_ = lo0111 & new_n5083_;
  assign new_n13106_ = ~new_n13099_ & ~new_n13104_;
  assign new_n13107_ = ~new_n13105_ & new_n13106_;
  assign new_n13108_ = new_n5070_ & ~new_n13107_;
  assign new_n13109_ = new_n13089_ & new_n13092_;
  assign new_n13110_ = new_n13098_ & new_n13109_;
  assign new_n13111_ = ~new_n13108_ & new_n13110_;
  assign new_n13112_ = ~new_n5105_ & new_n13010_;
  assign new_n13113_ = new_n13111_ & ~new_n13112_;
  assign new_n13114_ = new_n3815_ & new_n13036_;
  assign new_n13115_ = new_n4088_ & new_n13012_;
  assign new_n13116_ = ~new_n13114_ & ~new_n13115_;
  assign new_n13117_ = new_n3820_ & new_n13010_;
  assign new_n13118_ = new_n3870_ & new_n13037_;
  assign new_n13119_ = ~new_n13117_ & ~new_n13118_;
  assign new_n13120_ = ~new_n4069_ & new_n13012_;
  assign new_n13121_ = new_n13119_ & ~new_n13120_;
  assign new_n13122_ = new_n13081_ & new_n13113_;
  assign new_n13123_ = new_n13116_ & new_n13122_;
  assign li0111 = ~new_n13121_ | ~new_n13123_;
  assign li0112 = lo0124 | lo0468;
  assign new_n13126_ = ~lo0113 & ~new_n6044_;
  assign new_n13127_ = lo0113 & new_n6044_;
  assign new_n13128_ = ~new_n13126_ & ~new_n13127_;
  assign new_n13129_ = new_n6028_ & new_n13128_;
  assign new_n13130_ = lo0113 & ~new_n6028_;
  assign new_n13131_ = ~new_n13129_ & ~new_n13130_;
  assign li0113 = new_n11966_ & ~new_n13131_;
  assign new_n13133_ = new_n3658_ & new_n6030_;
  assign new_n13134_ = ~lo0114 & ~new_n13133_;
  assign new_n13135_ = lo0114 & new_n13133_;
  assign new_n13136_ = ~new_n13134_ & ~new_n13135_;
  assign new_n13137_ = new_n6028_ & new_n13136_;
  assign new_n13138_ = lo0114 & ~new_n6028_;
  assign new_n13139_ = ~new_n13137_ & ~new_n13138_;
  assign li0114 = new_n11966_ & ~new_n13139_;
  assign new_n13141_ = ~lo0115 & ~new_n6929_;
  assign new_n13142_ = lo0115 & new_n6929_;
  assign new_n13143_ = ~new_n13141_ & ~new_n13142_;
  assign new_n13144_ = new_n6028_ & new_n13143_;
  assign new_n13145_ = lo0115 & ~new_n6028_;
  assign new_n13146_ = ~new_n13144_ & ~new_n13145_;
  assign li0115 = new_n11966_ & ~new_n13146_;
  assign new_n13148_ = ~lo0116 & ~new_n6085_;
  assign new_n13149_ = lo0116 & new_n6085_;
  assign new_n13150_ = ~new_n13148_ & ~new_n13149_;
  assign new_n13151_ = new_n6028_ & new_n13150_;
  assign new_n13152_ = lo0116 & ~new_n6028_;
  assign new_n13153_ = ~new_n13151_ & ~new_n13152_;
  assign li0116 = new_n11966_ & ~new_n13153_;
  assign new_n13155_ = new_n3801_ & new_n3850_;
  assign new_n13156_ = new_n3917_ & new_n13155_;
  assign new_n13157_ = ~new_n3922_ & new_n3943_;
  assign new_n13158_ = new_n3756_ & new_n13157_;
  assign new_n13159_ = new_n3880_ & new_n13158_;
  assign new_n13160_ = new_n4026_ & new_n13156_;
  assign new_n13161_ = new_n13159_ & new_n13160_;
  assign li0117 = ~new_n3729_ | ~new_n13161_;
  assign new_n13163_ = ~new_n4543_ & ~new_n5252_;
  assign new_n13164_ = ~new_n4364_ & ~new_n5252_;
  assign new_n13165_ = lo0185 & ~new_n3522_;
  assign new_n13166_ = lo0150 & ~lo0185;
  assign new_n13167_ = ~new_n13165_ & ~new_n13166_;
  assign new_n13168_ = new_n4543_ & new_n13167_;
  assign new_n13169_ = ~new_n9853_ & ~new_n9862_;
  assign new_n13170_ = ~new_n13168_ & ~new_n13169_;
  assign new_n13171_ = new_n13168_ & new_n13169_;
  assign new_n13172_ = ~new_n13170_ & ~new_n13171_;
  assign new_n13173_ = new_n5252_ & ~new_n13172_;
  assign new_n13174_ = ~new_n5297_ & new_n13173_;
  assign new_n13175_ = lo0143 & ~new_n3522_;
  assign new_n13176_ = ~lo0143 & lo0165;
  assign new_n13177_ = ~new_n13175_ & ~new_n13176_;
  assign new_n13178_ = new_n4543_ & new_n13177_;
  assign new_n13179_ = new_n5268_ & new_n5280_;
  assign new_n13180_ = ~lo0118 & new_n9840_;
  assign new_n13181_ = lo0118 & ~new_n9840_;
  assign new_n13182_ = ~new_n13180_ & ~new_n13181_;
  assign new_n13183_ = ~new_n5276_ & ~new_n13182_;
  assign new_n13184_ = lo0118 & new_n13182_;
  assign new_n13185_ = ~new_n13183_ & ~new_n13184_;
  assign new_n13186_ = ~new_n5268_ & ~new_n13178_;
  assign new_n13187_ = new_n13179_ & ~new_n13185_;
  assign new_n13188_ = ~new_n13186_ & ~new_n13187_;
  assign new_n13189_ = ~new_n5259_ & new_n5297_;
  assign new_n13190_ = ~new_n13168_ & new_n13189_;
  assign new_n13191_ = new_n9834_ & ~new_n13188_;
  assign new_n13192_ = new_n5297_ & new_n13191_;
  assign new_n13193_ = ~new_n13190_ & ~new_n13192_;
  assign new_n13194_ = new_n5252_ & ~new_n13193_;
  assign new_n13195_ = ~new_n13163_ & ~new_n13164_;
  assign new_n13196_ = ~new_n13174_ & new_n13195_;
  assign new_n13197_ = ~new_n13194_ & new_n13196_;
  assign new_n13198_ = ~new_n4250_ & new_n4543_;
  assign new_n13199_ = ~new_n5313_ & ~new_n13198_;
  assign new_n13200_ = new_n5313_ & ~new_n13197_;
  assign new_n13201_ = ~new_n13199_ & ~new_n13200_;
  assign new_n13202_ = ~new_n5245_ & ~new_n5302_;
  assign new_n13203_ = new_n5245_ & ~new_n13201_;
  assign li0118 = new_n13202_ | new_n13203_;
  assign new_n13205_ = ~new_n3799_ & ~new_n3979_;
  assign new_n13206_ = ~new_n4655_ & ~new_n11250_;
  assign new_n13207_ = ~new_n10563_ & new_n13206_;
  assign new_n13208_ = new_n4475_ & ~new_n13207_;
  assign new_n13209_ = new_n4527_ & new_n13208_;
  assign new_n13210_ = ~new_n4560_ & ~new_n13209_;
  assign new_n13211_ = ~new_n4007_ & new_n13210_;
  assign new_n13212_ = ~new_n11125_ & new_n13211_;
  assign new_n13213_ = ~new_n9554_ & new_n13212_;
  assign new_n13214_ = new_n13205_ & new_n13213_;
  assign new_n13215_ = ~new_n3699_ & ~new_n4050_;
  assign new_n13216_ = ~new_n3936_ & new_n13214_;
  assign new_n13217_ = new_n13215_ & new_n13216_;
  assign li0131 = new_n3862_ | ~new_n13217_;
  assign new_n13219_ = lo0128 & ~lo0228;
  assign new_n13220_ = ~lo0128 & li0131;
  assign li0119 = new_n13219_ | new_n13220_;
  assign new_n13222_ = ~lo0031 & ~lo0080;
  assign new_n13223_ = lo0818 & new_n13222_;
  assign new_n13224_ = ~lo0982 & new_n5051_;
  assign new_n13225_ = new_n3673_ & new_n13224_;
  assign new_n13226_ = ~lo0951 & new_n13225_;
  assign li0818 = new_n13223_ | new_n13226_;
  assign new_n13228_ = pi004 & li0818;
  assign new_n13229_ = ~lo0120 & ~new_n13228_;
  assign li0120 = ~li0122 & ~new_n13229_;
  assign new_n13231_ = new_n3612_ & new_n4427_;
  assign new_n13232_ = ~new_n3612_ & new_n3940_;
  assign new_n13233_ = ~new_n13231_ & ~new_n13232_;
  assign new_n13234_ = new_n3799_ & ~new_n3979_;
  assign new_n13235_ = ~lo0024 & new_n3979_;
  assign new_n13236_ = ~new_n13234_ & ~new_n13235_;
  assign new_n13237_ = ~new_n4543_ & ~new_n13236_;
  assign new_n13238_ = lo0087 & ~new_n12845_;
  assign new_n13239_ = ~new_n9853_ & new_n13238_;
  assign new_n13240_ = lo0051 & ~new_n4543_;
  assign new_n13241_ = lo0051 & ~new_n3653_;
  assign new_n13242_ = ~new_n13240_ & ~new_n13241_;
  assign new_n13243_ = ~lo0125 & ~lo0133;
  assign new_n13244_ = ~lo0121 & new_n13243_;
  assign new_n13245_ = lo0121 & ~new_n13243_;
  assign new_n13246_ = ~new_n13244_ & ~new_n13245_;
  assign new_n13247_ = ~lo0126 & ~lo0132;
  assign new_n13248_ = new_n13244_ & new_n13247_;
  assign new_n13249_ = ~lo0130 & new_n13248_;
  assign new_n13250_ = ~lo0136 & new_n13249_;
  assign new_n13251_ = ~lo0134 & ~lo0135;
  assign new_n13252_ = new_n13250_ & new_n13251_;
  assign new_n13253_ = ~new_n13246_ & ~new_n13252_;
  assign new_n13254_ = ~lo0084 & new_n3567_;
  assign new_n13255_ = ~lo0068 & new_n13254_;
  assign new_n13256_ = ~new_n5323_ & ~new_n13255_;
  assign new_n13257_ = new_n13253_ & new_n13255_;
  assign new_n13258_ = ~new_n13256_ & ~new_n13257_;
  assign new_n13259_ = ~lo0051 & ~lo0087;
  assign new_n13260_ = ~new_n13258_ & new_n13259_;
  assign new_n13261_ = ~lo0087 & ~new_n13242_;
  assign new_n13262_ = ~new_n13260_ & ~new_n13261_;
  assign new_n13263_ = ~new_n12845_ & ~new_n13262_;
  assign new_n13264_ = ~new_n13239_ & ~new_n13263_;
  assign new_n13265_ = new_n12845_ & new_n13236_;
  assign new_n13266_ = ~new_n4557_ & new_n13265_;
  assign new_n13267_ = new_n13236_ & ~new_n13264_;
  assign new_n13268_ = ~new_n13266_ & ~new_n13267_;
  assign new_n13269_ = ~new_n9878_ & ~new_n13236_;
  assign new_n13270_ = new_n13233_ & ~new_n13237_;
  assign new_n13271_ = new_n13268_ & new_n13270_;
  assign new_n13272_ = ~new_n13269_ & new_n13271_;
  assign new_n13273_ = new_n3612_ & new_n4428_;
  assign new_n13274_ = ~new_n13272_ & new_n13273_;
  assign new_n13275_ = ~new_n4548_ & new_n13272_;
  assign li0121 = new_n13274_ | new_n13275_;
  assign new_n13277_ = lo0068 & ~lo0081;
  assign new_n13278_ = ~lo0048 & new_n13277_;
  assign new_n13279_ = ~lo0083 & new_n3842_;
  assign new_n13280_ = ~lo0067 & ~lo0085;
  assign new_n13281_ = ~lo0069 & ~lo0071;
  assign new_n13282_ = ~lo0087 & ~lo0109;
  assign new_n13283_ = ~lo0077 & new_n13282_;
  assign new_n13284_ = ~lo0103 & new_n13283_;
  assign new_n13285_ = ~lo0072 & new_n13284_;
  assign new_n13286_ = ~lo0086 & new_n13285_;
  assign new_n13287_ = ~lo0036 & ~lo0110;
  assign new_n13288_ = new_n3544_ & new_n13287_;
  assign new_n13289_ = ~lo0073 & new_n13288_;
  assign new_n13290_ = ~lo0091 & new_n13289_;
  assign new_n13291_ = ~lo0090 & new_n3553_;
  assign new_n13292_ = ~lo0047 & new_n13291_;
  assign new_n13293_ = new_n13290_ & new_n13292_;
  assign new_n13294_ = ~lo0111 & new_n13293_;
  assign new_n13295_ = new_n13286_ & new_n13294_;
  assign new_n13296_ = new_n13281_ & new_n13295_;
  assign new_n13297_ = new_n13280_ & new_n13296_;
  assign new_n13298_ = new_n13279_ & new_n13297_;
  assign new_n13299_ = ~lo0066 & new_n13298_;
  assign new_n13300_ = lo0081 & new_n13299_;
  assign new_n13301_ = lo0067 & new_n13296_;
  assign new_n13302_ = ~lo0085 & new_n13301_;
  assign new_n13303_ = new_n3553_ & new_n3851_;
  assign new_n13304_ = lo0073 & new_n13291_;
  assign new_n13305_ = ~new_n13303_ & ~new_n13304_;
  assign new_n13306_ = new_n4170_ & ~new_n13305_;
  assign new_n13307_ = ~lo0111 & new_n3549_;
  assign new_n13308_ = lo0111 & new_n13293_;
  assign new_n13309_ = new_n13306_ & new_n13307_;
  assign new_n13310_ = ~new_n13308_ & ~new_n13309_;
  assign new_n13311_ = ~lo0072 & ~new_n13294_;
  assign new_n13312_ = new_n13294_ & new_n13310_;
  assign new_n13313_ = ~new_n13311_ & ~new_n13312_;
  assign new_n13314_ = new_n4166_ & new_n13313_;
  assign new_n13315_ = new_n4165_ & new_n4175_;
  assign new_n13316_ = lo0071 & ~lo0085;
  assign new_n13317_ = ~lo0069 & new_n13316_;
  assign new_n13318_ = lo0069 & new_n4175_;
  assign new_n13319_ = ~new_n13317_ & ~new_n13318_;
  assign new_n13320_ = lo0085 & new_n13281_;
  assign new_n13321_ = new_n13295_ & ~new_n13319_;
  assign new_n13322_ = new_n13295_ & new_n13320_;
  assign new_n13323_ = ~new_n13321_ & ~new_n13322_;
  assign new_n13324_ = new_n13314_ & new_n13315_;
  assign new_n13325_ = new_n13323_ & ~new_n13324_;
  assign new_n13326_ = ~lo0067 & ~new_n13325_;
  assign new_n13327_ = ~new_n13302_ & ~new_n13326_;
  assign new_n13328_ = ~lo0083 & ~new_n13327_;
  assign new_n13329_ = lo0083 & new_n13297_;
  assign new_n13330_ = ~new_n13328_ & ~new_n13329_;
  assign new_n13331_ = new_n3837_ & new_n13297_;
  assign new_n13332_ = ~lo0083 & new_n13331_;
  assign new_n13333_ = new_n3557_ & new_n13332_;
  assign new_n13334_ = new_n3559_ & ~new_n13330_;
  assign new_n13335_ = ~new_n13333_ & ~new_n13334_;
  assign new_n13336_ = lo0066 & new_n13298_;
  assign new_n13337_ = new_n13335_ & ~new_n13336_;
  assign new_n13338_ = ~lo0081 & ~new_n13337_;
  assign new_n13339_ = ~new_n13300_ & ~new_n13338_;
  assign new_n13340_ = ~lo0048 & ~lo0068;
  assign new_n13341_ = ~new_n13339_ & new_n13340_;
  assign new_n13342_ = new_n13278_ & new_n13299_;
  assign new_n13343_ = ~new_n13341_ & ~new_n13342_;
  assign new_n13344_ = ~lo0059 & ~lo0062;
  assign new_n13345_ = ~li0893 & new_n13344_;
  assign new_n13346_ = ~lo0065 & new_n4149_;
  assign new_n13347_ = new_n4153_ & new_n13346_;
  assign new_n13348_ = new_n4189_ & new_n13347_;
  assign new_n13349_ = ~lo0057 & new_n13348_;
  assign new_n13350_ = new_n13345_ & new_n13349_;
  assign new_n13351_ = ~new_n13343_ & new_n13350_;
  assign new_n13352_ = new_n4194_ & new_n13351_;
  assign new_n13353_ = ~lo0074 & ~lo0094;
  assign new_n13354_ = new_n3527_ & new_n13353_;
  assign new_n13355_ = ~lo0096 & ~lo0097;
  assign new_n13356_ = new_n13354_ & new_n13355_;
  assign new_n13357_ = new_n5297_ & new_n13356_;
  assign new_n13358_ = new_n13352_ & new_n13357_;
  assign new_n13359_ = ~lo0045 & ~lo0055;
  assign new_n13360_ = new_n4158_ & new_n13359_;
  assign new_n13361_ = ~lo0038 & ~lo0053;
  assign new_n13362_ = new_n3573_ & new_n13361_;
  assign new_n13363_ = new_n13360_ & new_n13362_;
  assign new_n13364_ = ~lo0056 & new_n13363_;
  assign new_n13365_ = new_n13358_ & new_n13364_;
  assign new_n13366_ = lo0039 & lo0110;
  assign new_n13367_ = ~lo0039 & ~lo0110;
  assign new_n13368_ = ~new_n13366_ & ~new_n13367_;
  assign new_n13369_ = ~new_n13365_ & ~new_n13368_;
  assign new_n13370_ = ~new_n5230_ & new_n13368_;
  assign new_n13371_ = lo0039 & ~lo0110;
  assign new_n13372_ = new_n13370_ & ~new_n13371_;
  assign new_n13373_ = ~new_n4529_ & ~new_n9359_;
  assign new_n13374_ = new_n4475_ & ~new_n13373_;
  assign new_n13375_ = new_n4526_ & new_n13374_;
  assign new_n13376_ = new_n4524_ & new_n13375_;
  assign new_n13377_ = ~lo0039 & lo0110;
  assign new_n13378_ = ~new_n13376_ & ~new_n13377_;
  assign new_n13379_ = new_n13368_ & new_n13378_;
  assign new_n13380_ = ~new_n13372_ & ~new_n13379_;
  assign new_n13381_ = new_n13370_ & ~new_n13376_;
  assign new_n13382_ = ~new_n13369_ & new_n13380_;
  assign li0124 = new_n13381_ | ~new_n13382_;
  assign new_n13384_ = lo0051 & ~new_n4279_;
  assign new_n13385_ = ~new_n13240_ & ~new_n13384_;
  assign new_n13386_ = lo0125 & lo0133;
  assign new_n13387_ = ~new_n13243_ & ~new_n13386_;
  assign new_n13388_ = new_n13255_ & ~new_n13387_;
  assign new_n13389_ = ~new_n5253_ & ~new_n13255_;
  assign new_n13390_ = ~new_n13252_ & new_n13388_;
  assign new_n13391_ = ~new_n13389_ & ~new_n13390_;
  assign new_n13392_ = new_n13259_ & ~new_n13391_;
  assign new_n13393_ = ~lo0087 & ~new_n13385_;
  assign new_n13394_ = ~new_n13392_ & ~new_n13393_;
  assign new_n13395_ = ~new_n12845_ & ~new_n13394_;
  assign new_n13396_ = ~new_n5346_ & new_n13238_;
  assign new_n13397_ = ~new_n13395_ & ~new_n13396_;
  assign new_n13398_ = new_n13236_ & ~new_n13397_;
  assign new_n13399_ = ~new_n4544_ & new_n13265_;
  assign new_n13400_ = ~new_n13398_ & ~new_n13399_;
  assign new_n13401_ = ~new_n5371_ & ~new_n13236_;
  assign new_n13402_ = new_n13400_ & ~new_n13401_;
  assign new_n13403_ = ~new_n13237_ & new_n13402_;
  assign new_n13404_ = new_n13233_ & ~new_n13273_;
  assign new_n13405_ = ~new_n4557_ & new_n13273_;
  assign new_n13406_ = ~new_n13403_ & new_n13404_;
  assign li0125 = new_n13405_ | new_n13406_;
  assign new_n13408_ = ~new_n13168_ & new_n13238_;
  assign new_n13409_ = lo0051 & ~new_n3525_;
  assign new_n13410_ = ~new_n13240_ & ~new_n13409_;
  assign new_n13411_ = ~lo0126 & new_n13244_;
  assign new_n13412_ = lo0126 & ~new_n13244_;
  assign new_n13413_ = ~new_n13411_ & ~new_n13412_;
  assign new_n13414_ = ~new_n13252_ & ~new_n13413_;
  assign new_n13415_ = lo0126 & new_n13252_;
  assign new_n13416_ = ~new_n13414_ & ~new_n13415_;
  assign new_n13417_ = ~new_n6037_ & ~new_n13255_;
  assign new_n13418_ = new_n13255_ & ~new_n13416_;
  assign new_n13419_ = ~new_n13417_ & ~new_n13418_;
  assign new_n13420_ = new_n13259_ & ~new_n13419_;
  assign new_n13421_ = ~lo0087 & ~new_n13410_;
  assign new_n13422_ = ~new_n13420_ & ~new_n13421_;
  assign new_n13423_ = ~new_n12845_ & ~new_n13422_;
  assign new_n13424_ = ~new_n13408_ & ~new_n13423_;
  assign new_n13425_ = ~new_n4548_ & new_n13265_;
  assign new_n13426_ = new_n13236_ & ~new_n13424_;
  assign new_n13427_ = ~new_n13425_ & ~new_n13426_;
  assign new_n13428_ = ~new_n5302_ & new_n13233_;
  assign new_n13429_ = ~new_n13236_ & new_n13428_;
  assign new_n13430_ = new_n13233_ & ~new_n13427_;
  assign new_n13431_ = ~new_n13429_ & ~new_n13430_;
  assign new_n13432_ = new_n13273_ & ~new_n13431_;
  assign new_n13433_ = ~new_n4553_ & new_n13431_;
  assign li0126 = new_n13432_ | new_n13433_;
  assign new_n13435_ = new_n4647_ & ~new_n5131_;
  assign new_n13436_ = lo0250 & new_n13435_;
  assign new_n13437_ = ~li0583 & ~new_n13436_;
  assign new_n13438_ = lo0127 & li0583;
  assign new_n13439_ = ~new_n13437_ & ~new_n13438_;
  assign new_n13440_ = new_n3755_ & new_n4024_;
  assign new_n13441_ = new_n3849_ & ~new_n3879_;
  assign new_n13442_ = ~new_n4068_ & new_n4492_;
  assign new_n13443_ = ~new_n3815_ & new_n13442_;
  assign new_n13444_ = new_n3872_ & new_n13443_;
  assign new_n13445_ = new_n13441_ & new_n13444_;
  assign new_n13446_ = ~new_n3618_ & ~new_n4088_;
  assign new_n13447_ = ~new_n3804_ & new_n13445_;
  assign new_n13448_ = new_n13446_ & new_n13447_;
  assign new_n13449_ = new_n3892_ & new_n3904_;
  assign new_n13450_ = new_n3800_ & new_n13449_;
  assign new_n13451_ = new_n3915_ & new_n13450_;
  assign new_n13452_ = new_n4043_ & new_n13451_;
  assign new_n13453_ = ~new_n3769_ & ~new_n4050_;
  assign new_n13454_ = ~new_n3777_ & ~new_n3780_;
  assign new_n13455_ = new_n13453_ & new_n13454_;
  assign new_n13456_ = new_n13452_ & new_n13455_;
  assign new_n13457_ = new_n4013_ & ~new_n4133_;
  assign new_n13458_ = new_n13456_ & new_n13457_;
  assign new_n13459_ = new_n6389_ & new_n13458_;
  assign new_n13460_ = new_n13448_ & new_n13459_;
  assign new_n13461_ = ~new_n3625_ & new_n5201_;
  assign new_n13462_ = ~new_n3723_ & new_n13461_;
  assign new_n13463_ = ~new_n3699_ & ~new_n3705_;
  assign new_n13464_ = new_n3941_ & new_n13463_;
  assign new_n13465_ = new_n4116_ & new_n13464_;
  assign new_n13466_ = new_n13462_ & new_n13465_;
  assign new_n13467_ = new_n13440_ & new_n13460_;
  assign new_n13468_ = new_n3613_ & new_n13467_;
  assign new_n13469_ = new_n13466_ & new_n13468_;
  assign new_n13470_ = ~new_n3705_ & ~new_n13439_;
  assign new_n13471_ = new_n13439_ & ~new_n13469_;
  assign new_n13472_ = ~new_n13470_ & ~new_n13471_;
  assign li0127 = lo0129 & ~new_n13472_;
  assign new_n13474_ = new_n4647_ & new_n6021_;
  assign new_n13475_ = lo0129 & new_n13474_;
  assign new_n13476_ = ~lo0129 & ~li0583;
  assign new_n13477_ = ~new_n13475_ & ~new_n13476_;
  assign new_n13478_ = ~new_n3699_ & new_n4050_;
  assign new_n13479_ = ~new_n13477_ & new_n13478_;
  assign new_n13480_ = new_n3699_ & new_n4050_;
  assign new_n13481_ = ~new_n13215_ & ~new_n13480_;
  assign new_n13482_ = ~new_n3723_ & new_n5201_;
  assign new_n13483_ = ~new_n3927_ & new_n13482_;
  assign new_n13484_ = new_n13465_ & new_n13483_;
  assign new_n13485_ = new_n13460_ & new_n13484_;
  assign new_n13486_ = new_n3613_ & new_n13485_;
  assign new_n13487_ = new_n13440_ & new_n13486_;
  assign new_n13488_ = ~lo0250 & ~li0583;
  assign new_n13489_ = lo0129 & lo0250;
  assign new_n13490_ = ~new_n13488_ & ~new_n13489_;
  assign new_n13491_ = new_n3699_ & ~new_n13490_;
  assign new_n13492_ = ~new_n13481_ & ~new_n13487_;
  assign new_n13493_ = ~new_n4050_ & new_n13491_;
  assign new_n13494_ = ~new_n13492_ & ~new_n13493_;
  assign li0129 = new_n13479_ | ~new_n13494_;
  assign new_n13496_ = ~new_n5346_ & new_n13273_;
  assign new_n13497_ = ~new_n12845_ & ~new_n13273_;
  assign new_n13498_ = lo0130 & ~new_n13248_;
  assign new_n13499_ = ~new_n13249_ & ~new_n13498_;
  assign new_n13500_ = ~new_n13252_ & ~new_n13499_;
  assign new_n13501_ = new_n13255_ & new_n13500_;
  assign new_n13502_ = ~lo0051 & ~new_n5261_;
  assign new_n13503_ = ~new_n13255_ & new_n13502_;
  assign new_n13504_ = ~lo0051 & new_n13501_;
  assign new_n13505_ = ~new_n13503_ & ~new_n13504_;
  assign new_n13506_ = ~lo0087 & new_n13505_;
  assign new_n13507_ = lo0087 & new_n5336_;
  assign new_n13508_ = ~new_n13506_ & ~new_n13507_;
  assign new_n13509_ = new_n13233_ & new_n13497_;
  assign new_n13510_ = new_n13236_ & new_n13509_;
  assign new_n13511_ = new_n13508_ & new_n13510_;
  assign li0130 = new_n13496_ | new_n13511_;
  assign new_n13513_ = new_n13236_ & new_n13404_;
  assign new_n13514_ = lo0051 & ~new_n13198_;
  assign new_n13515_ = ~lo0121 & ~lo0126;
  assign new_n13516_ = new_n13243_ & new_n13515_;
  assign new_n13517_ = ~lo0132 & new_n13516_;
  assign new_n13518_ = lo0132 & ~new_n13516_;
  assign new_n13519_ = ~new_n13517_ & ~new_n13518_;
  assign new_n13520_ = lo0132 & ~new_n13252_;
  assign new_n13521_ = ~lo0132 & ~new_n13519_;
  assign new_n13522_ = ~new_n13520_ & ~new_n13521_;
  assign new_n13523_ = ~lo0051 & new_n13255_;
  assign new_n13524_ = ~new_n4364_ & ~new_n13255_;
  assign new_n13525_ = ~new_n4543_ & ~new_n13255_;
  assign new_n13526_ = ~new_n13524_ & ~new_n13525_;
  assign new_n13527_ = ~lo0051 & ~new_n13526_;
  assign new_n13528_ = ~new_n13522_ & new_n13523_;
  assign new_n13529_ = ~new_n13527_ & ~new_n13528_;
  assign new_n13530_ = ~new_n13514_ & new_n13529_;
  assign new_n13531_ = ~lo0087 & ~new_n12845_;
  assign new_n13532_ = ~new_n4553_ & new_n12845_;
  assign new_n13533_ = ~new_n5265_ & new_n13238_;
  assign new_n13534_ = ~new_n13532_ & ~new_n13533_;
  assign new_n13535_ = ~new_n13530_ & new_n13531_;
  assign new_n13536_ = new_n13534_ & ~new_n13535_;
  assign new_n13537_ = ~new_n5293_ & new_n13273_;
  assign new_n13538_ = new_n13513_ & ~new_n13536_;
  assign li0132 = new_n13537_ | new_n13538_;
  assign new_n13540_ = ~new_n12845_ & new_n13236_;
  assign new_n13541_ = ~lo0133 & new_n13252_;
  assign new_n13542_ = lo0133 & ~new_n13252_;
  assign new_n13543_ = ~new_n13541_ & ~new_n13542_;
  assign new_n13544_ = new_n13523_ & ~new_n13543_;
  assign new_n13545_ = ~lo0087 & ~new_n13544_;
  assign new_n13546_ = lo0087 & ~new_n5293_;
  assign new_n13547_ = ~new_n13545_ & ~new_n13546_;
  assign new_n13548_ = new_n13540_ & ~new_n13547_;
  assign new_n13549_ = ~new_n4235_ & ~new_n13236_;
  assign new_n13550_ = ~new_n13548_ & ~new_n13549_;
  assign new_n13551_ = ~new_n13237_ & new_n13550_;
  assign new_n13552_ = new_n13404_ & ~new_n13551_;
  assign new_n13553_ = ~new_n4544_ & new_n13273_;
  assign li0133 = new_n13552_ | new_n13553_;
  assign new_n13555_ = ~lo0135 & ~lo0136;
  assign new_n13556_ = ~lo0130 & ~lo0132;
  assign new_n13557_ = new_n13516_ & new_n13555_;
  assign new_n13558_ = new_n13556_ & new_n13557_;
  assign new_n13559_ = lo0134 & ~new_n13558_;
  assign new_n13560_ = ~lo0134 & new_n13558_;
  assign new_n13561_ = ~new_n13559_ & ~new_n13560_;
  assign new_n13562_ = ~new_n13252_ & ~new_n13561_;
  assign new_n13563_ = lo0134 & new_n13252_;
  assign new_n13564_ = ~new_n13562_ & ~new_n13563_;
  assign new_n13565_ = new_n13255_ & ~new_n13564_;
  assign new_n13566_ = ~new_n4296_ & ~new_n13255_;
  assign new_n13567_ = ~new_n13565_ & ~new_n13566_;
  assign new_n13568_ = ~new_n13525_ & new_n13567_;
  assign new_n13569_ = new_n13236_ & ~new_n13568_;
  assign new_n13570_ = ~new_n12845_ & new_n13259_;
  assign new_n13571_ = new_n13569_ & new_n13570_;
  assign new_n13572_ = new_n13404_ & new_n13571_;
  assign new_n13573_ = ~new_n5265_ & new_n13273_;
  assign li0134 = new_n13572_ | new_n13573_;
  assign new_n13575_ = ~lo0130 & new_n13244_;
  assign new_n13576_ = ~lo0136 & new_n13247_;
  assign new_n13577_ = new_n13575_ & new_n13576_;
  assign new_n13578_ = ~lo0135 & new_n13577_;
  assign new_n13579_ = lo0135 & ~new_n13577_;
  assign new_n13580_ = ~new_n13578_ & ~new_n13579_;
  assign new_n13581_ = ~new_n13252_ & ~new_n13580_;
  assign new_n13582_ = lo0135 & new_n13252_;
  assign new_n13583_ = ~new_n13581_ & ~new_n13582_;
  assign new_n13584_ = new_n13255_ & ~new_n13583_;
  assign new_n13585_ = ~new_n4313_ & ~new_n13255_;
  assign new_n13586_ = ~new_n13584_ & ~new_n13585_;
  assign new_n13587_ = ~new_n13525_ & new_n13586_;
  assign new_n13588_ = new_n13236_ & ~new_n13587_;
  assign new_n13589_ = new_n13570_ & new_n13588_;
  assign new_n13590_ = new_n13404_ & new_n13589_;
  assign new_n13591_ = ~new_n13168_ & new_n13273_;
  assign li0135 = new_n13590_ | new_n13591_;
  assign new_n13593_ = new_n13515_ & new_n13556_;
  assign new_n13594_ = new_n13243_ & new_n13593_;
  assign new_n13595_ = lo0136 & ~new_n13594_;
  assign new_n13596_ = ~lo0136 & new_n13594_;
  assign new_n13597_ = ~new_n13595_ & ~new_n13596_;
  assign new_n13598_ = lo0136 & ~new_n13252_;
  assign new_n13599_ = ~lo0136 & ~new_n13597_;
  assign new_n13600_ = ~new_n13598_ & ~new_n13599_;
  assign new_n13601_ = ~new_n13255_ & ~new_n13600_;
  assign new_n13602_ = ~new_n5324_ & new_n13600_;
  assign new_n13603_ = ~new_n13601_ & ~new_n13602_;
  assign new_n13604_ = ~new_n13273_ & ~new_n13603_;
  assign new_n13605_ = new_n13236_ & new_n13604_;
  assign new_n13606_ = new_n13233_ & new_n13605_;
  assign new_n13607_ = ~new_n9853_ & new_n13273_;
  assign new_n13608_ = new_n13570_ & new_n13606_;
  assign li0136 = new_n13607_ | new_n13608_;
  assign new_n13610_ = new_n4053_ & new_n6103_;
  assign new_n13611_ = ~lo0039 & lo0137;
  assign li0137 = new_n13610_ | new_n13611_;
  assign new_n13613_ = ~new_n5252_ & ~new_n5324_;
  assign new_n13614_ = new_n5280_ & new_n5297_;
  assign new_n13615_ = new_n9834_ & new_n13614_;
  assign new_n13616_ = lo0138 & ~new_n5272_;
  assign new_n13617_ = ~new_n5273_ & ~new_n13616_;
  assign new_n13618_ = new_n5276_ & ~new_n13617_;
  assign new_n13619_ = lo0138 & ~new_n5276_;
  assign new_n13620_ = ~new_n13618_ & ~new_n13619_;
  assign new_n13621_ = new_n5252_ & new_n13615_;
  assign new_n13622_ = new_n5268_ & new_n13621_;
  assign new_n13623_ = ~new_n13620_ & new_n13622_;
  assign new_n13624_ = new_n5245_ & new_n5313_;
  assign new_n13625_ = ~new_n13613_ & ~new_n13623_;
  assign li0138 = new_n13624_ & ~new_n13625_;
  assign new_n13627_ = ~new_n5252_ & ~new_n5261_;
  assign new_n13628_ = new_n5269_ & new_n5325_;
  assign new_n13629_ = ~lo0139 & new_n13628_;
  assign new_n13630_ = lo0139 & ~new_n13628_;
  assign new_n13631_ = ~new_n13629_ & ~new_n13630_;
  assign new_n13632_ = new_n5276_ & ~new_n13631_;
  assign new_n13633_ = lo0139 & ~new_n5276_;
  assign new_n13634_ = ~new_n13632_ & ~new_n13633_;
  assign new_n13635_ = new_n13622_ & ~new_n13634_;
  assign new_n13636_ = ~new_n13627_ & ~new_n13635_;
  assign li0139 = new_n13624_ & ~new_n13636_;
  assign new_n13638_ = ~lo0120 & li0583;
  assign new_n13639_ = lo0120 & new_n4219_;
  assign new_n13640_ = new_n5076_ & ~new_n13639_;
  assign new_n13641_ = ~new_n13638_ & ~new_n13640_;
  assign new_n13642_ = new_n4475_ & new_n13641_;
  assign new_n13643_ = lo0120 & ~new_n4475_;
  assign new_n13644_ = ~new_n13642_ & ~new_n13643_;
  assign new_n13645_ = ~lo0979 & new_n4526_;
  assign new_n13646_ = new_n13644_ & new_n13645_;
  assign new_n13647_ = new_n4653_ & ~new_n13646_;
  assign new_n13648_ = new_n4023_ & new_n5222_;
  assign new_n13649_ = new_n4091_ & new_n13648_;
  assign new_n13650_ = ~li0793 & new_n13649_;
  assign new_n13651_ = lo0120 & lo0287;
  assign new_n13652_ = new_n3612_ & new_n13651_;
  assign new_n13653_ = ~new_n4018_ & ~new_n13652_;
  assign new_n13654_ = ~new_n3773_ & new_n13653_;
  assign new_n13655_ = ~new_n13650_ & new_n13654_;
  assign new_n13656_ = ~new_n9215_ & new_n13655_;
  assign new_n13657_ = lo0841 & ~li0583;
  assign new_n13658_ = new_n3867_ & new_n13657_;
  assign new_n13659_ = ~new_n3996_ & ~new_n13658_;
  assign new_n13660_ = lo0252 & ~new_n13659_;
  assign new_n13661_ = ~new_n3618_ & ~new_n3879_;
  assign new_n13662_ = lo0252 & new_n5211_;
  assign new_n13663_ = new_n4004_ & new_n13662_;
  assign new_n13664_ = new_n13661_ & ~new_n13663_;
  assign new_n13665_ = ~new_n13647_ & new_n13656_;
  assign new_n13666_ = ~new_n13660_ & new_n13665_;
  assign li0230 = ~new_n13664_ | ~new_n13666_;
  assign new_n13668_ = new_n3673_ & li0230;
  assign new_n13669_ = lo0832 & new_n3673_;
  assign new_n13670_ = ~new_n13668_ & ~new_n13669_;
  assign new_n13671_ = lo0738 & ~new_n13670_;
  assign new_n13672_ = lo0609 & lo0785;
  assign new_n13673_ = pi066 & lo0785;
  assign new_n13674_ = ~new_n13672_ & ~new_n13673_;
  assign new_n13675_ = lo0609 & new_n13672_;
  assign new_n13676_ = ~new_n13674_ & ~new_n13675_;
  assign new_n13677_ = ~lo0785 & ~new_n13673_;
  assign new_n13678_ = pi064 & lo0778;
  assign new_n13679_ = lo0778 & new_n13678_;
  assign new_n13680_ = lo0608 & new_n13679_;
  assign new_n13681_ = ~lo0608 & ~new_n13678_;
  assign new_n13682_ = ~new_n13680_ & ~new_n13681_;
  assign new_n13683_ = ~lo0778 & ~new_n13678_;
  assign new_n13684_ = new_n13682_ & ~new_n13683_;
  assign new_n13685_ = ~new_n13676_ & ~new_n13677_;
  assign new_n13686_ = ~new_n13684_ & ~new_n13685_;
  assign new_n13687_ = pi065 & lo0781;
  assign new_n13688_ = ~lo0781 & ~new_n13687_;
  assign new_n13689_ = ~lo0618 & ~new_n13687_;
  assign new_n13690_ = lo0618 & new_n13687_;
  assign new_n13691_ = lo0781 & new_n13690_;
  assign new_n13692_ = ~new_n13688_ & ~new_n13689_;
  assign new_n13693_ = ~new_n13691_ & new_n13692_;
  assign new_n13694_ = lo0629 & lo0792;
  assign new_n13695_ = pi067 & lo0792;
  assign new_n13696_ = ~new_n13694_ & ~new_n13695_;
  assign new_n13697_ = lo0629 & new_n13694_;
  assign new_n13698_ = ~new_n13696_ & ~new_n13697_;
  assign new_n13699_ = ~lo0792 & ~new_n13695_;
  assign new_n13700_ = pi071 & lo0790;
  assign new_n13701_ = ~lo0790 & ~new_n13700_;
  assign new_n13702_ = ~lo0644 & ~new_n13700_;
  assign new_n13703_ = lo0644 & lo0790;
  assign new_n13704_ = new_n13700_ & new_n13703_;
  assign new_n13705_ = ~new_n13701_ & ~new_n13702_;
  assign new_n13706_ = ~new_n13704_ & new_n13705_;
  assign new_n13707_ = lo0603 & ~new_n13706_;
  assign new_n13708_ = ~new_n13698_ & ~new_n13699_;
  assign new_n13709_ = new_n13707_ & ~new_n13708_;
  assign new_n13710_ = lo0630 & lo0787;
  assign new_n13711_ = pi068 & lo0787;
  assign new_n13712_ = ~new_n13710_ & ~new_n13711_;
  assign new_n13713_ = lo0630 & new_n13710_;
  assign new_n13714_ = ~new_n13712_ & ~new_n13713_;
  assign new_n13715_ = ~lo0787 & ~new_n13711_;
  assign new_n13716_ = pi070 & lo0789;
  assign new_n13717_ = lo0619 & new_n13716_;
  assign new_n13718_ = lo0789 & new_n13717_;
  assign new_n13719_ = ~lo0619 & ~new_n13716_;
  assign new_n13720_ = ~new_n13718_ & ~new_n13719_;
  assign new_n13721_ = ~lo0789 & ~new_n13716_;
  assign new_n13722_ = pi069 & lo0788;
  assign new_n13723_ = ~lo0788 & ~new_n13722_;
  assign new_n13724_ = ~lo0626 & ~new_n13722_;
  assign new_n13725_ = lo0626 & lo0788;
  assign new_n13726_ = new_n13722_ & new_n13725_;
  assign new_n13727_ = ~new_n13723_ & ~new_n13724_;
  assign new_n13728_ = ~new_n13726_ & new_n13727_;
  assign new_n13729_ = new_n13720_ & ~new_n13721_;
  assign new_n13730_ = ~new_n13728_ & ~new_n13729_;
  assign new_n13731_ = ~new_n13714_ & ~new_n13715_;
  assign new_n13732_ = new_n13730_ & ~new_n13731_;
  assign new_n13733_ = new_n13686_ & ~new_n13693_;
  assign new_n13734_ = new_n13709_ & new_n13733_;
  assign new_n13735_ = new_n13732_ & new_n13734_;
  assign new_n13736_ = pi002 & lo0621;
  assign new_n13737_ = new_n13735_ & ~new_n13736_;
  assign new_n13738_ = lo0628 & lo0792;
  assign new_n13739_ = ~new_n13695_ & ~new_n13738_;
  assign new_n13740_ = lo0628 & new_n13738_;
  assign new_n13741_ = ~new_n13739_ & ~new_n13740_;
  assign new_n13742_ = lo0627 & lo0781;
  assign new_n13743_ = ~new_n13687_ & ~new_n13742_;
  assign new_n13744_ = lo0627 & new_n13742_;
  assign new_n13745_ = ~new_n13743_ & ~new_n13744_;
  assign new_n13746_ = ~new_n13699_ & ~new_n13741_;
  assign new_n13747_ = ~new_n13688_ & ~new_n13745_;
  assign new_n13748_ = ~new_n13746_ & ~new_n13747_;
  assign new_n13749_ = ~lo0660 & ~new_n13673_;
  assign new_n13750_ = lo0660 & new_n13673_;
  assign new_n13751_ = lo0785 & new_n13750_;
  assign new_n13752_ = ~new_n13677_ & ~new_n13749_;
  assign new_n13753_ = ~new_n13751_ & new_n13752_;
  assign new_n13754_ = lo0715 & lo0790;
  assign new_n13755_ = ~new_n13700_ & ~new_n13754_;
  assign new_n13756_ = lo0715 & new_n13754_;
  assign new_n13757_ = ~new_n13755_ & ~new_n13756_;
  assign new_n13758_ = lo0625 & new_n13679_;
  assign new_n13759_ = ~lo0625 & ~new_n13678_;
  assign new_n13760_ = ~new_n13758_ & ~new_n13759_;
  assign new_n13761_ = ~new_n13683_ & new_n13760_;
  assign new_n13762_ = lo0680 & ~new_n13761_;
  assign new_n13763_ = ~new_n13701_ & ~new_n13757_;
  assign new_n13764_ = new_n13762_ & ~new_n13763_;
  assign new_n13765_ = lo0641 & lo0788;
  assign new_n13766_ = ~new_n13722_ & ~new_n13765_;
  assign new_n13767_ = lo0641 & new_n13765_;
  assign new_n13768_ = ~new_n13766_ & ~new_n13767_;
  assign new_n13769_ = lo0648 & new_n13716_;
  assign new_n13770_ = lo0789 & new_n13769_;
  assign new_n13771_ = ~lo0648 & ~new_n13716_;
  assign new_n13772_ = ~new_n13770_ & ~new_n13771_;
  assign new_n13773_ = ~lo0647 & ~new_n13711_;
  assign new_n13774_ = lo0647 & new_n13711_;
  assign new_n13775_ = lo0787 & new_n13774_;
  assign new_n13776_ = ~new_n13715_ & ~new_n13773_;
  assign new_n13777_ = ~new_n13775_ & new_n13776_;
  assign new_n13778_ = ~new_n13721_ & new_n13772_;
  assign new_n13779_ = ~new_n13777_ & ~new_n13778_;
  assign new_n13780_ = ~new_n13723_ & ~new_n13768_;
  assign new_n13781_ = new_n13779_ & ~new_n13780_;
  assign new_n13782_ = new_n13748_ & ~new_n13753_;
  assign new_n13783_ = new_n13764_ & new_n13782_;
  assign new_n13784_ = new_n13781_ & new_n13783_;
  assign new_n13785_ = pi002 & lo0665;
  assign new_n13786_ = new_n13784_ & ~new_n13785_;
  assign new_n13787_ = ~new_n13737_ & new_n13786_;
  assign new_n13788_ = lo0761 & new_n13737_;
  assign new_n13789_ = ~new_n13670_ & new_n13788_;
  assign new_n13790_ = new_n13671_ & new_n13787_;
  assign new_n13791_ = ~new_n13789_ & ~new_n13790_;
  assign new_n13792_ = lo0140 & new_n13670_;
  assign li0140 = ~new_n13791_ | new_n13792_;
  assign new_n13794_ = lo0706 & ~new_n13670_;
  assign new_n13795_ = lo0749 & new_n13737_;
  assign new_n13796_ = ~new_n13670_ & new_n13795_;
  assign new_n13797_ = new_n13787_ & new_n13794_;
  assign new_n13798_ = ~new_n13796_ & ~new_n13797_;
  assign new_n13799_ = lo0141 & new_n13670_;
  assign li0141 = ~new_n13798_ | new_n13799_;
  assign new_n13801_ = lo0735 & ~new_n13670_;
  assign new_n13802_ = lo0743 & new_n13737_;
  assign new_n13803_ = ~new_n13670_ & new_n13802_;
  assign new_n13804_ = new_n13787_ & new_n13801_;
  assign new_n13805_ = ~new_n13803_ & ~new_n13804_;
  assign new_n13806_ = lo0142 & new_n13670_;
  assign li0142 = ~new_n13805_ | new_n13806_;
  assign new_n13808_ = lo0687 & ~new_n13670_;
  assign new_n13809_ = lo0774 & new_n13737_;
  assign new_n13810_ = ~new_n13670_ & new_n13809_;
  assign new_n13811_ = new_n13787_ & new_n13808_;
  assign new_n13812_ = ~new_n13810_ & ~new_n13811_;
  assign new_n13813_ = lo0143 & new_n13670_;
  assign li0143 = ~new_n13812_ | new_n13813_;
  assign new_n13815_ = lo0736 & ~new_n13670_;
  assign new_n13816_ = lo0758 & new_n13737_;
  assign new_n13817_ = ~new_n13670_ & new_n13816_;
  assign new_n13818_ = new_n13787_ & new_n13815_;
  assign new_n13819_ = ~new_n13817_ & ~new_n13818_;
  assign new_n13820_ = lo0144 & new_n13670_;
  assign li0144 = ~new_n13819_ | new_n13820_;
  assign new_n13822_ = lo0698 & ~new_n13670_;
  assign new_n13823_ = lo0767 & new_n13737_;
  assign new_n13824_ = ~new_n13670_ & new_n13823_;
  assign new_n13825_ = new_n13787_ & new_n13822_;
  assign new_n13826_ = ~new_n13824_ & ~new_n13825_;
  assign new_n13827_ = lo0145 & new_n13670_;
  assign li0145 = ~new_n13826_ | new_n13827_;
  assign new_n13829_ = lo0907 & ~lo0947;
  assign new_n13830_ = lo0743 & lo0947;
  assign new_n13831_ = ~new_n13670_ & new_n13830_;
  assign new_n13832_ = new_n13801_ & new_n13829_;
  assign new_n13833_ = ~new_n13831_ & ~new_n13832_;
  assign new_n13834_ = lo0146 & new_n13670_;
  assign li0146 = ~new_n13833_ | new_n13834_;
  assign new_n13836_ = lo0726 & ~new_n13670_;
  assign new_n13837_ = lo0770 & lo0947;
  assign new_n13838_ = ~new_n13670_ & new_n13837_;
  assign new_n13839_ = new_n13829_ & new_n13836_;
  assign new_n13840_ = ~new_n13838_ & ~new_n13839_;
  assign new_n13841_ = lo0147 & new_n13670_;
  assign li0147 = ~new_n13840_ | new_n13841_;
  assign new_n13843_ = lo0749 & lo0947;
  assign new_n13844_ = ~new_n13670_ & new_n13843_;
  assign new_n13845_ = new_n13794_ & new_n13829_;
  assign new_n13846_ = ~new_n13844_ & ~new_n13845_;
  assign new_n13847_ = lo0148 & new_n13670_;
  assign li0148 = ~new_n13846_ | new_n13847_;
  assign new_n13849_ = lo0725 & ~new_n13670_;
  assign new_n13850_ = lo0755 & lo0947;
  assign new_n13851_ = ~new_n13670_ & new_n13850_;
  assign new_n13852_ = new_n13829_ & new_n13849_;
  assign new_n13853_ = ~new_n13851_ & ~new_n13852_;
  assign new_n13854_ = lo0149 & new_n13670_;
  assign li0149 = ~new_n13853_ | new_n13854_;
  assign new_n13856_ = lo0701 & ~new_n13670_;
  assign new_n13857_ = lo0751 & lo0947;
  assign new_n13858_ = ~new_n13670_ & new_n13857_;
  assign new_n13859_ = new_n13829_ & new_n13856_;
  assign new_n13860_ = ~new_n13858_ & ~new_n13859_;
  assign new_n13861_ = lo0150 & new_n13670_;
  assign li0150 = ~new_n13860_ | new_n13861_;
  assign new_n13863_ = lo0723 & ~new_n13670_;
  assign new_n13864_ = lo0745 & lo0947;
  assign new_n13865_ = ~new_n13670_ & new_n13864_;
  assign new_n13866_ = new_n13829_ & new_n13863_;
  assign new_n13867_ = ~new_n13865_ & ~new_n13866_;
  assign new_n13868_ = lo0151 & new_n13670_;
  assign li0151 = ~new_n13867_ | new_n13868_;
  assign new_n13870_ = lo0696 & ~new_n13670_;
  assign new_n13871_ = lo0759 & lo0947;
  assign new_n13872_ = ~new_n13670_ & new_n13871_;
  assign new_n13873_ = new_n13829_ & new_n13870_;
  assign new_n13874_ = ~new_n13872_ & ~new_n13873_;
  assign new_n13875_ = lo0152 & new_n13670_;
  assign li0152 = ~new_n13874_ | new_n13875_;
  assign new_n13877_ = lo0700 & ~new_n13670_;
  assign new_n13878_ = lo0766 & lo0947;
  assign new_n13879_ = ~new_n13670_ & new_n13878_;
  assign new_n13880_ = new_n13829_ & new_n13877_;
  assign new_n13881_ = ~new_n13879_ & ~new_n13880_;
  assign new_n13882_ = lo0153 & new_n13670_;
  assign li0153 = ~new_n13881_ | new_n13882_;
  assign new_n13884_ = lo0704 & ~new_n13670_;
  assign new_n13885_ = lo0742 & lo0947;
  assign new_n13886_ = ~new_n13670_ & new_n13885_;
  assign new_n13887_ = new_n13829_ & new_n13884_;
  assign new_n13888_ = ~new_n13886_ & ~new_n13887_;
  assign new_n13889_ = lo0154 & new_n13670_;
  assign li0154 = ~new_n13888_ | new_n13889_;
  assign new_n13891_ = lo0686 & ~new_n13670_;
  assign new_n13892_ = lo0757 & lo0947;
  assign new_n13893_ = ~new_n13670_ & new_n13892_;
  assign new_n13894_ = new_n13829_ & new_n13891_;
  assign new_n13895_ = ~new_n13893_ & ~new_n13894_;
  assign new_n13896_ = lo0155 & new_n13670_;
  assign li0155 = ~new_n13895_ | new_n13896_;
  assign new_n13898_ = lo0724 & ~new_n13670_;
  assign new_n13899_ = lo0741 & lo0947;
  assign new_n13900_ = ~new_n13670_ & new_n13899_;
  assign new_n13901_ = new_n13829_ & new_n13898_;
  assign new_n13902_ = ~new_n13900_ & ~new_n13901_;
  assign new_n13903_ = lo0156 & new_n13670_;
  assign li0156 = ~new_n13902_ | new_n13903_;
  assign new_n13905_ = lo0688 & ~new_n13670_;
  assign new_n13906_ = lo0760 & lo0947;
  assign new_n13907_ = ~new_n13670_ & new_n13906_;
  assign new_n13908_ = new_n13829_ & new_n13905_;
  assign new_n13909_ = ~new_n13907_ & ~new_n13908_;
  assign new_n13910_ = lo0157 & new_n13670_;
  assign li0157 = ~new_n13909_ | new_n13910_;
  assign new_n13912_ = lo0702 & ~new_n13670_;
  assign new_n13913_ = lo0753 & lo0947;
  assign new_n13914_ = ~new_n13670_ & new_n13913_;
  assign new_n13915_ = new_n13829_ & new_n13912_;
  assign new_n13916_ = ~new_n13914_ & ~new_n13915_;
  assign new_n13917_ = lo0158 & new_n13670_;
  assign li0158 = ~new_n13916_ | new_n13917_;
  assign new_n13919_ = lo0709 & ~new_n13670_;
  assign new_n13920_ = lo0754 & lo0947;
  assign new_n13921_ = ~new_n13670_ & new_n13920_;
  assign new_n13922_ = new_n13829_ & new_n13919_;
  assign new_n13923_ = ~new_n13921_ & ~new_n13922_;
  assign new_n13924_ = lo0159 & new_n13670_;
  assign li0159 = ~new_n13923_ | new_n13924_;
  assign new_n13926_ = lo0734 & ~new_n13670_;
  assign new_n13927_ = lo0756 & lo0947;
  assign new_n13928_ = ~new_n13670_ & new_n13927_;
  assign new_n13929_ = new_n13829_ & new_n13926_;
  assign new_n13930_ = ~new_n13928_ & ~new_n13929_;
  assign new_n13931_ = lo0160 & new_n13670_;
  assign li0160 = ~new_n13930_ | new_n13931_;
  assign new_n13933_ = lo0758 & lo0947;
  assign new_n13934_ = ~new_n13670_ & new_n13933_;
  assign new_n13935_ = new_n13815_ & new_n13829_;
  assign new_n13936_ = ~new_n13934_ & ~new_n13935_;
  assign new_n13937_ = lo0161 & new_n13670_;
  assign li0161 = ~new_n13936_ | new_n13937_;
  assign new_n13939_ = lo0761 & lo0947;
  assign new_n13940_ = ~new_n13670_ & new_n13939_;
  assign new_n13941_ = new_n13671_ & new_n13829_;
  assign new_n13942_ = ~new_n13940_ & ~new_n13941_;
  assign new_n13943_ = lo0162 & new_n13670_;
  assign li0162 = ~new_n13942_ | new_n13943_;
  assign new_n13945_ = lo0737 & ~new_n13670_;
  assign new_n13946_ = lo0777 & lo0947;
  assign new_n13947_ = ~new_n13670_ & new_n13946_;
  assign new_n13948_ = new_n13829_ & new_n13945_;
  assign new_n13949_ = ~new_n13947_ & ~new_n13948_;
  assign new_n13950_ = lo0163 & new_n13670_;
  assign li0163 = ~new_n13949_ | new_n13950_;
  assign new_n13952_ = lo0703 & ~new_n13670_;
  assign new_n13953_ = lo0752 & lo0947;
  assign new_n13954_ = ~new_n13670_ & new_n13953_;
  assign new_n13955_ = new_n13829_ & new_n13952_;
  assign new_n13956_ = ~new_n13954_ & ~new_n13955_;
  assign new_n13957_ = lo0164 & new_n13670_;
  assign li0164 = ~new_n13956_ | new_n13957_;
  assign new_n13959_ = lo0774 & lo0947;
  assign new_n13960_ = ~new_n13670_ & new_n13959_;
  assign new_n13961_ = new_n13808_ & new_n13829_;
  assign new_n13962_ = ~new_n13960_ & ~new_n13961_;
  assign new_n13963_ = lo0165 & new_n13670_;
  assign li0165 = ~new_n13962_ | new_n13963_;
  assign new_n13965_ = lo0727 & ~new_n13670_;
  assign new_n13966_ = lo0772 & lo0947;
  assign new_n13967_ = ~new_n13670_ & new_n13966_;
  assign new_n13968_ = new_n13829_ & new_n13965_;
  assign new_n13969_ = ~new_n13967_ & ~new_n13968_;
  assign new_n13970_ = lo0166 & new_n13670_;
  assign li0166 = ~new_n13969_ | new_n13970_;
  assign new_n13972_ = lo0705 & ~new_n13670_;
  assign new_n13973_ = lo0768 & lo0947;
  assign new_n13974_ = ~new_n13670_ & new_n13973_;
  assign new_n13975_ = new_n13829_ & new_n13972_;
  assign new_n13976_ = ~new_n13974_ & ~new_n13975_;
  assign new_n13977_ = lo0167 & new_n13670_;
  assign li0167 = ~new_n13976_ | new_n13977_;
  assign new_n13979_ = lo0699 & ~new_n13670_;
  assign new_n13980_ = lo0763 & lo0947;
  assign new_n13981_ = ~new_n13670_ & new_n13980_;
  assign new_n13982_ = new_n13829_ & new_n13979_;
  assign new_n13983_ = ~new_n13981_ & ~new_n13982_;
  assign new_n13984_ = lo0168 & new_n13670_;
  assign li0168 = ~new_n13983_ | new_n13984_;
  assign new_n13986_ = lo0729 & ~new_n13670_;
  assign new_n13987_ = lo0746 & lo0947;
  assign new_n13988_ = ~new_n13670_ & new_n13987_;
  assign new_n13989_ = new_n13829_ & new_n13986_;
  assign new_n13990_ = ~new_n13988_ & ~new_n13989_;
  assign new_n13991_ = lo0169 & new_n13670_;
  assign li0169 = ~new_n13990_ | new_n13991_;
  assign new_n13993_ = lo0730 & ~new_n13670_;
  assign new_n13994_ = lo0748 & lo0947;
  assign new_n13995_ = ~new_n13670_ & new_n13994_;
  assign new_n13996_ = new_n13829_ & new_n13993_;
  assign new_n13997_ = ~new_n13995_ & ~new_n13996_;
  assign new_n13998_ = lo0170 & new_n13670_;
  assign li0170 = ~new_n13997_ | new_n13998_;
  assign new_n14000_ = lo0691 & ~new_n13670_;
  assign new_n14001_ = lo0764 & lo0947;
  assign new_n14002_ = ~new_n13670_ & new_n14001_;
  assign new_n14003_ = new_n13829_ & new_n14000_;
  assign new_n14004_ = ~new_n14002_ & ~new_n14003_;
  assign new_n14005_ = lo0171 & new_n13670_;
  assign li0171 = ~new_n14004_ | new_n14005_;
  assign new_n14007_ = lo0690 & ~new_n13670_;
  assign new_n14008_ = lo0739 & lo0947;
  assign new_n14009_ = ~new_n13670_ & new_n14008_;
  assign new_n14010_ = new_n13829_ & new_n14007_;
  assign new_n14011_ = ~new_n14009_ & ~new_n14010_;
  assign new_n14012_ = lo0172 & new_n13670_;
  assign li0172 = ~new_n14011_ | new_n14012_;
  assign new_n14014_ = lo0745 & new_n13737_;
  assign new_n14015_ = ~new_n13670_ & new_n14014_;
  assign new_n14016_ = new_n13787_ & new_n13863_;
  assign new_n14017_ = ~new_n14015_ & ~new_n14016_;
  assign new_n14018_ = lo0173 & new_n13670_;
  assign li0173 = ~new_n14017_ | new_n14018_;
  assign new_n14020_ = lo0759 & new_n13737_;
  assign new_n14021_ = ~new_n13670_ & new_n14020_;
  assign new_n14022_ = new_n13787_ & new_n13870_;
  assign new_n14023_ = ~new_n14021_ & ~new_n14022_;
  assign new_n14024_ = lo0174 & new_n13670_;
  assign li0174 = ~new_n14023_ | new_n14024_;
  assign new_n14026_ = lo0766 & new_n13737_;
  assign new_n14027_ = ~new_n13670_ & new_n14026_;
  assign new_n14028_ = new_n13787_ & new_n13877_;
  assign new_n14029_ = ~new_n14027_ & ~new_n14028_;
  assign new_n14030_ = lo0175 & new_n13670_;
  assign li0175 = ~new_n14029_ | new_n14030_;
  assign new_n14032_ = lo0742 & new_n13737_;
  assign new_n14033_ = ~new_n13670_ & new_n14032_;
  assign new_n14034_ = new_n13787_ & new_n13884_;
  assign new_n14035_ = ~new_n14033_ & ~new_n14034_;
  assign new_n14036_ = lo0176 & new_n13670_;
  assign li0176 = ~new_n14035_ | new_n14036_;
  assign new_n14038_ = lo0757 & new_n13737_;
  assign new_n14039_ = ~new_n13670_ & new_n14038_;
  assign new_n14040_ = new_n13787_ & new_n13891_;
  assign new_n14041_ = ~new_n14039_ & ~new_n14040_;
  assign new_n14042_ = lo0177 & new_n13670_;
  assign li0177 = ~new_n14041_ | new_n14042_;
  assign new_n14044_ = lo0760 & new_n13737_;
  assign new_n14045_ = ~new_n13670_ & new_n14044_;
  assign new_n14046_ = new_n13787_ & new_n13905_;
  assign new_n14047_ = ~new_n14045_ & ~new_n14046_;
  assign new_n14048_ = lo0178 & new_n13670_;
  assign li0178 = ~new_n14047_ | new_n14048_;
  assign new_n14050_ = lo0741 & new_n13737_;
  assign new_n14051_ = ~new_n13670_ & new_n14050_;
  assign new_n14052_ = new_n13787_ & new_n13898_;
  assign new_n14053_ = ~new_n14051_ & ~new_n14052_;
  assign new_n14054_ = lo0179 & new_n13670_;
  assign li0179 = ~new_n14053_ | new_n14054_;
  assign new_n14056_ = lo0753 & new_n13737_;
  assign new_n14057_ = ~new_n13670_ & new_n14056_;
  assign new_n14058_ = new_n13787_ & new_n13912_;
  assign new_n14059_ = ~new_n14057_ & ~new_n14058_;
  assign new_n14060_ = lo0180 & new_n13670_;
  assign li0180 = ~new_n14059_ | new_n14060_;
  assign new_n14062_ = lo0754 & new_n13737_;
  assign new_n14063_ = ~new_n13670_ & new_n14062_;
  assign new_n14064_ = new_n13787_ & new_n13919_;
  assign new_n14065_ = ~new_n14063_ & ~new_n14064_;
  assign new_n14066_ = lo0181 & new_n13670_;
  assign li0181 = ~new_n14065_ | new_n14066_;
  assign new_n14068_ = lo0756 & new_n13737_;
  assign new_n14069_ = ~new_n13670_ & new_n14068_;
  assign new_n14070_ = new_n13787_ & new_n13926_;
  assign new_n14071_ = ~new_n14069_ & ~new_n14070_;
  assign new_n14072_ = lo0182 & new_n13670_;
  assign li0182 = ~new_n14071_ | new_n14072_;
  assign new_n14074_ = lo0755 & new_n13737_;
  assign new_n14075_ = ~new_n13670_ & new_n14074_;
  assign new_n14076_ = new_n13787_ & new_n13849_;
  assign new_n14077_ = ~new_n14075_ & ~new_n14076_;
  assign new_n14078_ = lo0183 & new_n13670_;
  assign li0183 = ~new_n14077_ | new_n14078_;
  assign new_n14080_ = lo0777 & new_n13737_;
  assign new_n14081_ = ~new_n13670_ & new_n14080_;
  assign new_n14082_ = new_n13787_ & new_n13945_;
  assign new_n14083_ = ~new_n14081_ & ~new_n14082_;
  assign new_n14084_ = lo0184 & new_n13670_;
  assign li0184 = ~new_n14083_ | new_n14084_;
  assign new_n14086_ = lo0751 & new_n13737_;
  assign new_n14087_ = ~new_n13670_ & new_n14086_;
  assign new_n14088_ = new_n13787_ & new_n13856_;
  assign new_n14089_ = ~new_n14087_ & ~new_n14088_;
  assign new_n14090_ = lo0185 & new_n13670_;
  assign li0185 = ~new_n14089_ | new_n14090_;
  assign new_n14092_ = lo0752 & new_n13737_;
  assign new_n14093_ = ~new_n13670_ & new_n14092_;
  assign new_n14094_ = new_n13787_ & new_n13952_;
  assign new_n14095_ = ~new_n14093_ & ~new_n14094_;
  assign new_n14096_ = lo0186 & new_n13670_;
  assign li0186 = ~new_n14095_ | new_n14096_;
  assign new_n14098_ = lo0770 & new_n13737_;
  assign new_n14099_ = ~new_n13670_ & new_n14098_;
  assign new_n14100_ = new_n13787_ & new_n13836_;
  assign new_n14101_ = ~new_n14099_ & ~new_n14100_;
  assign new_n14102_ = lo0187 & new_n13670_;
  assign li0187 = ~new_n14101_ | new_n14102_;
  assign new_n14104_ = lo0768 & new_n13737_;
  assign new_n14105_ = ~new_n13670_ & new_n14104_;
  assign new_n14106_ = new_n13787_ & new_n13972_;
  assign new_n14107_ = ~new_n14105_ & ~new_n14106_;
  assign new_n14108_ = lo0188 & new_n13670_;
  assign li0188 = ~new_n14107_ | new_n14108_;
  assign new_n14110_ = lo0772 & new_n13737_;
  assign new_n14111_ = ~new_n13670_ & new_n14110_;
  assign new_n14112_ = new_n13787_ & new_n13965_;
  assign new_n14113_ = ~new_n14111_ & ~new_n14112_;
  assign new_n14114_ = lo0189 & new_n13670_;
  assign li0189 = ~new_n14113_ | new_n14114_;
  assign new_n14116_ = lo0763 & new_n13737_;
  assign new_n14117_ = ~new_n13670_ & new_n14116_;
  assign new_n14118_ = new_n13787_ & new_n13979_;
  assign new_n14119_ = ~new_n14117_ & ~new_n14118_;
  assign new_n14120_ = lo0190 & new_n13670_;
  assign li0190 = ~new_n14119_ | new_n14120_;
  assign new_n14122_ = lo0746 & new_n13737_;
  assign new_n14123_ = ~new_n13670_ & new_n14122_;
  assign new_n14124_ = new_n13787_ & new_n13986_;
  assign new_n14125_ = ~new_n14123_ & ~new_n14124_;
  assign new_n14126_ = lo0191 & new_n13670_;
  assign li0191 = ~new_n14125_ | new_n14126_;
  assign new_n14128_ = lo0764 & new_n13737_;
  assign new_n14129_ = ~new_n13670_ & new_n14128_;
  assign new_n14130_ = new_n13787_ & new_n14000_;
  assign new_n14131_ = ~new_n14129_ & ~new_n14130_;
  assign new_n14132_ = lo0192 & new_n13670_;
  assign li0192 = ~new_n14131_ | new_n14132_;
  assign new_n14134_ = lo0739 & new_n13737_;
  assign new_n14135_ = ~new_n13670_ & new_n14134_;
  assign new_n14136_ = new_n13787_ & new_n14007_;
  assign new_n14137_ = ~new_n14135_ & ~new_n14136_;
  assign new_n14138_ = lo0193 & new_n13670_;
  assign li0193 = ~new_n14137_ | new_n14138_;
  assign new_n14140_ = lo0748 & new_n13737_;
  assign new_n14141_ = ~new_n13670_ & new_n14140_;
  assign new_n14142_ = new_n13787_ & new_n13993_;
  assign new_n14143_ = ~new_n14141_ & ~new_n14142_;
  assign new_n14144_ = lo0194 & new_n13670_;
  assign li0194 = ~new_n14143_ | new_n14144_;
  assign new_n14146_ = ~lo0138 & ~lo0196;
  assign new_n14147_ = ~lo0139 & new_n9840_;
  assign new_n14148_ = ~lo0118 & new_n14147_;
  assign new_n14149_ = new_n14146_ & new_n14148_;
  assign new_n14150_ = ~lo0195 & ~new_n14149_;
  assign new_n14151_ = lo0195 & new_n14149_;
  assign new_n14152_ = ~new_n14150_ & ~new_n14151_;
  assign new_n14153_ = new_n5276_ & new_n14152_;
  assign new_n14154_ = lo0195 & ~new_n5276_;
  assign new_n14155_ = ~new_n14153_ & ~new_n14154_;
  assign new_n14156_ = new_n5268_ & ~new_n14155_;
  assign new_n14157_ = new_n5252_ & new_n14156_;
  assign new_n14158_ = new_n5280_ & new_n14157_;
  assign new_n14159_ = new_n9833_ & new_n14158_;
  assign new_n14160_ = new_n5259_ & new_n5297_;
  assign new_n14161_ = new_n14159_ & new_n14160_;
  assign new_n14162_ = ~new_n4296_ & ~new_n5252_;
  assign new_n14163_ = ~new_n14161_ & ~new_n14162_;
  assign new_n14164_ = ~new_n13163_ & new_n14163_;
  assign li0195 = new_n13624_ & ~new_n14164_;
  assign new_n14166_ = ~lo0139 & new_n5325_;
  assign new_n14167_ = ~lo0138 & new_n14166_;
  assign new_n14168_ = new_n5269_ & new_n14167_;
  assign new_n14169_ = ~lo0196 & ~new_n14168_;
  assign new_n14170_ = lo0196 & new_n14168_;
  assign new_n14171_ = ~new_n14169_ & ~new_n14170_;
  assign new_n14172_ = new_n5276_ & new_n14171_;
  assign new_n14173_ = lo0196 & ~new_n5276_;
  assign new_n14174_ = ~new_n14172_ & ~new_n14173_;
  assign new_n14175_ = new_n5268_ & ~new_n14174_;
  assign new_n14176_ = new_n5252_ & new_n14175_;
  assign new_n14177_ = new_n13615_ & new_n14176_;
  assign new_n14178_ = ~new_n4313_ & ~new_n5252_;
  assign new_n14179_ = ~new_n14177_ & ~new_n14178_;
  assign new_n14180_ = ~new_n13163_ & new_n14179_;
  assign li0196 = new_n13624_ & ~new_n14180_;
  assign new_n14182_ = lo0767 & lo0947;
  assign new_n14183_ = ~new_n13670_ & new_n14182_;
  assign new_n14184_ = new_n13822_ & new_n13829_;
  assign new_n14185_ = ~new_n14183_ & ~new_n14184_;
  assign new_n14186_ = lo0197 & new_n13670_;
  assign li0197 = ~new_n14185_ | new_n14186_;
  assign new_n14188_ = lo0198 & ~new_n13668_;
  assign new_n14189_ = lo0634 & new_n13668_;
  assign new_n14190_ = new_n13787_ & new_n14189_;
  assign new_n14191_ = new_n13668_ & new_n13737_;
  assign new_n14192_ = lo0633 & new_n14191_;
  assign new_n14193_ = ~new_n14188_ & ~new_n14190_;
  assign li0198 = new_n14192_ | ~new_n14193_;
  assign new_n14195_ = lo0199 & ~new_n13668_;
  assign new_n14196_ = lo0637 & new_n13668_;
  assign new_n14197_ = new_n13787_ & new_n14196_;
  assign new_n14198_ = lo0617 & new_n14191_;
  assign new_n14199_ = ~new_n14195_ & ~new_n14197_;
  assign li0199 = new_n14198_ | ~new_n14199_;
  assign new_n14201_ = lo0200 & ~new_n13668_;
  assign new_n14202_ = lo0643 & new_n13668_;
  assign new_n14203_ = new_n13787_ & new_n14202_;
  assign new_n14204_ = lo0606 & new_n14191_;
  assign new_n14205_ = ~new_n14201_ & ~new_n14203_;
  assign li0200 = new_n14204_ | ~new_n14205_;
  assign new_n14207_ = ~lo0032 & lo0070;
  assign new_n14208_ = ~lo0332 & new_n14207_;
  assign new_n14209_ = lo0032 & ~lo0070;
  assign new_n14210_ = new_n4534_ & new_n14209_;
  assign new_n14211_ = ~new_n14208_ & ~new_n14210_;
  assign new_n14212_ = new_n4460_ & ~new_n14211_;
  assign new_n14213_ = ~lo0233 & ~lo0237;
  assign new_n14214_ = new_n14212_ & new_n14213_;
  assign new_n14215_ = lo0201 & ~lo0332;
  assign new_n14216_ = ~new_n14214_ & new_n14215_;
  assign new_n14217_ = ~lo0053 & ~lo0106;
  assign new_n14218_ = new_n4168_ & new_n4184_;
  assign new_n14219_ = ~lo0088 & new_n14218_;
  assign new_n14220_ = new_n3549_ & new_n14219_;
  assign new_n14221_ = ~lo0092 & new_n14220_;
  assign new_n14222_ = ~lo0047 & new_n14221_;
  assign new_n14223_ = new_n3548_ & new_n14222_;
  assign new_n14224_ = ~lo0058 & new_n14223_;
  assign new_n14225_ = ~lo0103 & new_n4164_;
  assign new_n14226_ = new_n4171_ & new_n14225_;
  assign new_n14227_ = ~lo0087 & new_n14226_;
  assign new_n14228_ = new_n4163_ & new_n4175_;
  assign new_n14229_ = ~lo0107 & new_n14228_;
  assign new_n14230_ = new_n3559_ & new_n4178_;
  assign new_n14231_ = new_n3578_ & new_n3581_;
  assign new_n14232_ = ~lo0063 & new_n14231_;
  assign new_n14233_ = new_n4149_ & new_n14229_;
  assign new_n14234_ = new_n14230_ & new_n14233_;
  assign new_n14235_ = new_n14232_ & new_n14234_;
  assign new_n14236_ = new_n14227_ & new_n14235_;
  assign new_n14237_ = new_n4176_ & new_n14224_;
  assign new_n14238_ = new_n14236_ & new_n14237_;
  assign new_n14239_ = ~lo0060 & new_n14238_;
  assign new_n14240_ = new_n3781_ & new_n14238_;
  assign new_n14241_ = lo0059 & new_n14239_;
  assign new_n14242_ = ~new_n14240_ & ~new_n14241_;
  assign new_n14243_ = new_n3575_ & ~new_n14242_;
  assign new_n14244_ = new_n4154_ & new_n14239_;
  assign new_n14245_ = new_n13344_ & new_n14244_;
  assign new_n14246_ = ~lo0045 & lo0055;
  assign new_n14247_ = new_n14245_ & new_n14246_;
  assign new_n14248_ = ~lo0045 & new_n14243_;
  assign new_n14249_ = new_n3520_ & new_n14248_;
  assign new_n14250_ = ~new_n14247_ & ~new_n14249_;
  assign new_n14251_ = new_n13359_ & new_n14245_;
  assign new_n14252_ = lo0054 & ~new_n14250_;
  assign new_n14253_ = new_n14250_ & new_n14251_;
  assign new_n14254_ = ~new_n14252_ & ~new_n14253_;
  assign new_n14255_ = lo0053 & new_n3573_;
  assign new_n14256_ = new_n14217_ & ~new_n14254_;
  assign new_n14257_ = new_n14251_ & new_n14255_;
  assign new_n14258_ = ~new_n14256_ & ~new_n14257_;
  assign new_n14259_ = ~lo0070 & new_n4189_;
  assign new_n14260_ = ~lo0096 & new_n14259_;
  assign new_n14261_ = ~new_n14258_ & new_n14260_;
  assign new_n14262_ = new_n3536_ & new_n4182_;
  assign new_n14263_ = new_n14261_ & new_n14262_;
  assign new_n14264_ = new_n3535_ & new_n14263_;
  assign new_n14265_ = ~lo0108 & new_n3540_;
  assign new_n14266_ = ~lo0035 & new_n14265_;
  assign new_n14267_ = new_n14264_ & new_n14266_;
  assign new_n14268_ = new_n4186_ & new_n4195_;
  assign new_n14269_ = ~lo0070 & new_n14268_;
  assign new_n14270_ = new_n14267_ & new_n14269_;
  assign new_n14271_ = lo0070 & lo0332;
  assign new_n14272_ = ~new_n14270_ & ~new_n14271_;
  assign new_n14273_ = new_n4460_ & ~new_n14272_;
  assign new_n14274_ = new_n4460_ & new_n11654_;
  assign new_n14275_ = new_n14213_ & new_n14274_;
  assign new_n14276_ = new_n14216_ & ~new_n14273_;
  assign li0201 = new_n14275_ | new_n14276_;
  assign new_n14278_ = lo0233 & ~lo0237;
  assign new_n14279_ = new_n14212_ & new_n14278_;
  assign new_n14280_ = ~lo0332 & ~new_n14273_;
  assign new_n14281_ = ~new_n14279_ & new_n14280_;
  assign new_n14282_ = lo0202 & new_n14281_;
  assign new_n14283_ = new_n14274_ & new_n14278_;
  assign li0202 = new_n14282_ | new_n14283_;
  assign new_n14285_ = lo0233 & lo0237;
  assign new_n14286_ = new_n14212_ & new_n14285_;
  assign new_n14287_ = new_n14280_ & ~new_n14286_;
  assign new_n14288_ = lo0203 & new_n14287_;
  assign new_n14289_ = new_n14274_ & new_n14285_;
  assign li0203 = new_n14288_ | new_n14289_;
  assign new_n14291_ = ~new_n4469_ & ~new_n14211_;
  assign new_n14292_ = new_n14213_ & new_n14291_;
  assign new_n14293_ = lo0204 & ~lo0332;
  assign new_n14294_ = ~new_n14292_ & new_n14293_;
  assign new_n14295_ = ~new_n4469_ & ~new_n14272_;
  assign new_n14296_ = ~new_n4469_ & new_n11654_;
  assign new_n14297_ = new_n14213_ & new_n14296_;
  assign new_n14298_ = new_n14294_ & ~new_n14295_;
  assign li0204 = new_n14297_ | new_n14298_;
  assign new_n14300_ = new_n14278_ & new_n14291_;
  assign new_n14301_ = ~lo0332 & ~new_n14295_;
  assign new_n14302_ = ~new_n14300_ & new_n14301_;
  assign new_n14303_ = lo0205 & new_n14302_;
  assign new_n14304_ = new_n14278_ & new_n14296_;
  assign li0205 = new_n14303_ | new_n14304_;
  assign new_n14306_ = ~lo0233 & lo0237;
  assign new_n14307_ = new_n14291_ & new_n14306_;
  assign new_n14308_ = new_n14301_ & ~new_n14307_;
  assign new_n14309_ = lo0206 & new_n14308_;
  assign new_n14310_ = new_n14296_ & new_n14306_;
  assign li0206 = new_n14309_ | new_n14310_;
  assign new_n14312_ = lo0623 & new_n13668_;
  assign new_n14313_ = lo0710 & new_n13668_;
  assign new_n14314_ = new_n13737_ & new_n14312_;
  assign new_n14315_ = new_n13787_ & new_n14313_;
  assign new_n14316_ = ~new_n14314_ & ~new_n14315_;
  assign new_n14317_ = lo0207 & ~new_n13668_;
  assign li0207 = ~new_n14316_ | new_n14317_;
  assign new_n14319_ = lo0607 & new_n13668_;
  assign new_n14320_ = lo0638 & new_n13668_;
  assign new_n14321_ = new_n13737_ & new_n14319_;
  assign new_n14322_ = new_n13787_ & new_n14320_;
  assign new_n14323_ = ~new_n14321_ & ~new_n14322_;
  assign new_n14324_ = lo0208 & ~new_n13668_;
  assign li0208 = ~new_n14323_ | new_n14324_;
  assign new_n14326_ = lo0622 & new_n13668_;
  assign new_n14327_ = lo0639 & new_n13668_;
  assign new_n14328_ = new_n13737_ & new_n14326_;
  assign new_n14329_ = new_n13787_ & new_n14327_;
  assign new_n14330_ = ~new_n14328_ & ~new_n14329_;
  assign new_n14331_ = lo0209 & ~new_n13668_;
  assign li0209 = ~new_n14330_ | new_n14331_;
  assign new_n14333_ = lo0210 & ~new_n13668_;
  assign new_n14334_ = new_n13829_ & new_n14189_;
  assign new_n14335_ = lo0633 & new_n13668_;
  assign new_n14336_ = lo0947 & new_n14335_;
  assign new_n14337_ = ~new_n14333_ & ~new_n14334_;
  assign li0210 = new_n14336_ | ~new_n14337_;
  assign new_n14339_ = lo0211 & ~new_n13668_;
  assign new_n14340_ = new_n13829_ & new_n14202_;
  assign new_n14341_ = lo0606 & new_n13668_;
  assign new_n14342_ = lo0947 & new_n14341_;
  assign new_n14343_ = ~new_n14339_ & ~new_n14340_;
  assign li0211 = new_n14342_ | ~new_n14343_;
  assign new_n14345_ = lo0607 & lo0947;
  assign new_n14346_ = new_n13668_ & new_n14345_;
  assign new_n14347_ = new_n13829_ & new_n14320_;
  assign new_n14348_ = ~new_n14346_ & ~new_n14347_;
  assign new_n14349_ = lo0212 & ~new_n13668_;
  assign li0212 = ~new_n14348_ | new_n14349_;
  assign new_n14351_ = lo0622 & lo0947;
  assign new_n14352_ = new_n13668_ & new_n14351_;
  assign new_n14353_ = new_n13829_ & new_n14327_;
  assign new_n14354_ = ~new_n14352_ & ~new_n14353_;
  assign new_n14355_ = lo0213 & ~new_n13668_;
  assign li0213 = ~new_n14354_ | new_n14355_;
  assign new_n14357_ = lo0623 & lo0947;
  assign new_n14358_ = new_n13668_ & new_n14357_;
  assign new_n14359_ = new_n13829_ & new_n14313_;
  assign new_n14360_ = ~new_n14358_ & ~new_n14359_;
  assign new_n14361_ = lo0214 & ~new_n13668_;
  assign li0214 = ~new_n14360_ | new_n14361_;
  assign new_n14363_ = lo0215 & ~new_n13668_;
  assign new_n14364_ = lo0947 & new_n13668_;
  assign new_n14365_ = lo0642 & new_n14364_;
  assign new_n14366_ = lo0907 & new_n13668_;
  assign new_n14367_ = lo0681 & new_n14366_;
  assign new_n14368_ = ~lo0947 & new_n14367_;
  assign new_n14369_ = ~new_n14363_ & ~new_n14365_;
  assign li0215 = new_n14368_ | ~new_n14369_;
  assign new_n14371_ = lo0216 & ~new_n13668_;
  assign new_n14372_ = lo0614 & new_n14364_;
  assign new_n14373_ = lo0662 & new_n14366_;
  assign new_n14374_ = ~lo0947 & new_n14373_;
  assign new_n14375_ = ~new_n14371_ & ~new_n14372_;
  assign li0216 = new_n14374_ | ~new_n14375_;
  assign new_n14377_ = lo0612 & new_n13737_;
  assign new_n14378_ = lo0695 & new_n13787_;
  assign new_n14379_ = ~new_n14377_ & ~new_n14378_;
  assign new_n14380_ = new_n13668_ & ~new_n14379_;
  assign new_n14381_ = lo0217 & ~new_n13668_;
  assign li0217 = new_n14380_ | new_n14381_;
  assign new_n14383_ = new_n14285_ & new_n14291_;
  assign new_n14384_ = new_n14301_ & ~new_n14383_;
  assign new_n14385_ = lo0218 & new_n14384_;
  assign new_n14386_ = new_n14285_ & new_n14296_;
  assign li0218 = new_n14385_ | new_n14386_;
  assign new_n14388_ = lo0219 & ~new_n13668_;
  assign new_n14389_ = new_n13829_ & new_n14196_;
  assign new_n14390_ = lo0617 & new_n13668_;
  assign new_n14391_ = lo0947 & new_n14390_;
  assign new_n14392_ = ~new_n14388_ & ~new_n14389_;
  assign li0219 = new_n14391_ | ~new_n14392_;
  assign new_n14394_ = new_n14212_ & new_n14306_;
  assign new_n14395_ = new_n14280_ & ~new_n14394_;
  assign new_n14396_ = lo0220 & new_n14395_;
  assign new_n14397_ = new_n14274_ & new_n14306_;
  assign li0220 = new_n14396_ | new_n14397_;
  assign new_n14399_ = lo0221 & ~new_n13668_;
  assign new_n14400_ = lo0616 & new_n14364_;
  assign new_n14401_ = lo0661 & new_n14366_;
  assign new_n14402_ = ~lo0947 & new_n14401_;
  assign new_n14403_ = ~new_n14399_ & ~new_n14400_;
  assign li0221 = new_n14402_ | ~new_n14403_;
  assign new_n14405_ = lo0616 & new_n13737_;
  assign new_n14406_ = lo0661 & new_n13787_;
  assign new_n14407_ = ~new_n14405_ & ~new_n14406_;
  assign new_n14408_ = lo0222 & new_n13668_;
  assign new_n14409_ = ~lo0222 & ~new_n14407_;
  assign li0222 = new_n14408_ | new_n14409_;
  assign new_n14411_ = lo0642 & new_n13737_;
  assign new_n14412_ = lo0681 & new_n13787_;
  assign new_n14413_ = ~new_n14411_ & ~new_n14412_;
  assign new_n14414_ = lo0223 & new_n13668_;
  assign new_n14415_ = ~lo0223 & ~new_n14413_;
  assign li0223 = new_n14414_ | new_n14415_;
  assign new_n14417_ = lo0614 & new_n13737_;
  assign new_n14418_ = lo0662 & new_n13787_;
  assign new_n14419_ = ~new_n14417_ & ~new_n14418_;
  assign new_n14420_ = lo0224 & new_n13668_;
  assign new_n14421_ = ~lo0224 & ~new_n14419_;
  assign li0224 = new_n14420_ | new_n14421_;
  assign new_n14423_ = lo0479 & new_n4020_;
  assign new_n14424_ = new_n4500_ & new_n13456_;
  assign new_n14425_ = new_n13445_ & new_n14424_;
  assign new_n14426_ = ~new_n14423_ & new_n14425_;
  assign new_n14427_ = new_n4012_ & new_n14426_;
  assign new_n14428_ = new_n3756_ & new_n14427_;
  assign li0236 = ~new_n13484_ | ~new_n14428_;
  assign new_n14430_ = ~lo0228 & lo0231;
  assign new_n14431_ = ~lo0231 & li0236;
  assign li0226 = new_n14430_ | new_n14431_;
  assign new_n14433_ = new_n4427_ & new_n5250_;
  assign new_n14434_ = ~lo0287 & new_n4422_;
  assign new_n14435_ = new_n14433_ & new_n14434_;
  assign new_n14436_ = ~new_n3891_ & new_n3941_;
  assign new_n14437_ = ~new_n14435_ & new_n14436_;
  assign new_n14438_ = ~new_n3834_ & ~new_n3996_;
  assign new_n14439_ = ~new_n3996_ & ~new_n14435_;
  assign new_n14440_ = new_n3678_ & ~new_n4528_;
  assign new_n14441_ = new_n14439_ & new_n14440_;
  assign new_n14442_ = new_n14436_ & new_n14441_;
  assign new_n14443_ = ~new_n4528_ & new_n14438_;
  assign new_n14444_ = new_n14437_ & new_n14443_;
  assign new_n14445_ = ~new_n14442_ & ~new_n14444_;
  assign new_n14446_ = ~new_n3753_ & ~new_n3996_;
  assign new_n14447_ = ~new_n3753_ & ~new_n14435_;
  assign new_n14448_ = new_n14438_ & new_n14447_;
  assign new_n14449_ = new_n14436_ & new_n14448_;
  assign new_n14450_ = new_n3678_ & new_n14446_;
  assign new_n14451_ = new_n14437_ & new_n14450_;
  assign new_n14452_ = ~new_n14449_ & ~new_n14451_;
  assign new_n14453_ = new_n14445_ & new_n14452_;
  assign new_n14454_ = ~new_n6399_ & ~new_n14435_;
  assign new_n14455_ = new_n14446_ & new_n14454_;
  assign new_n14456_ = ~new_n3834_ & ~new_n3940_;
  assign new_n14457_ = ~new_n3936_ & new_n14456_;
  assign new_n14458_ = new_n3678_ & ~new_n6399_;
  assign new_n14459_ = new_n14447_ & new_n14458_;
  assign new_n14460_ = ~new_n3940_ & ~new_n3996_;
  assign new_n14461_ = ~new_n3936_ & new_n14460_;
  assign new_n14462_ = new_n14455_ & new_n14457_;
  assign new_n14463_ = new_n14459_ & new_n14461_;
  assign new_n14464_ = ~new_n14462_ & ~new_n14463_;
  assign new_n14465_ = ~new_n4528_ & ~new_n6399_;
  assign new_n14466_ = new_n14439_ & new_n14457_;
  assign new_n14467_ = new_n14465_ & new_n14466_;
  assign new_n14468_ = new_n14440_ & new_n14461_;
  assign new_n14469_ = new_n14454_ & new_n14468_;
  assign new_n14470_ = new_n14453_ & new_n14464_;
  assign new_n14471_ = ~new_n14467_ & new_n14470_;
  assign new_n14472_ = ~new_n14469_ & new_n14471_;
  assign new_n14473_ = ~new_n3612_ & ~new_n3936_;
  assign new_n14474_ = ~new_n3891_ & new_n14473_;
  assign new_n14475_ = ~new_n3996_ & new_n14474_;
  assign new_n14476_ = new_n14440_ & new_n14460_;
  assign new_n14477_ = new_n14474_ & new_n14476_;
  assign new_n14478_ = ~new_n4528_ & new_n14456_;
  assign new_n14479_ = new_n14475_ & new_n14478_;
  assign new_n14480_ = ~new_n14477_ & ~new_n14479_;
  assign new_n14481_ = new_n14472_ & new_n14480_;
  assign new_n14482_ = ~new_n3753_ & new_n14438_;
  assign new_n14483_ = ~new_n3612_ & new_n3941_;
  assign new_n14484_ = new_n14458_ & new_n14483_;
  assign new_n14485_ = new_n14446_ & new_n14484_;
  assign new_n14486_ = ~new_n6399_ & new_n14483_;
  assign new_n14487_ = new_n14482_ & new_n14486_;
  assign new_n14488_ = ~new_n14485_ & ~new_n14487_;
  assign new_n14489_ = new_n3678_ & new_n14460_;
  assign new_n14490_ = new_n14446_ & new_n14456_;
  assign new_n14491_ = new_n14474_ & new_n14490_;
  assign new_n14492_ = ~new_n3753_ & new_n14474_;
  assign new_n14493_ = new_n14489_ & new_n14492_;
  assign new_n14494_ = ~new_n14491_ & ~new_n14493_;
  assign new_n14495_ = new_n14488_ & new_n14494_;
  assign new_n14496_ = ~new_n3996_ & new_n14483_;
  assign new_n14497_ = ~new_n6399_ & new_n14440_;
  assign new_n14498_ = new_n14496_ & new_n14497_;
  assign new_n14499_ = new_n14465_ & new_n14483_;
  assign new_n14500_ = new_n14438_ & new_n14499_;
  assign new_n14501_ = new_n14481_ & new_n14495_;
  assign new_n14502_ = ~new_n14498_ & new_n14501_;
  assign li0227 = new_n14500_ | ~new_n14502_;
  assign new_n14504_ = ~lo0039 & lo0228;
  assign new_n14505_ = ~li0683 & ~new_n4666_;
  assign new_n14506_ = ~new_n3612_ & ~new_n3974_;
  assign new_n14507_ = ~new_n3810_ & ~new_n3974_;
  assign new_n14508_ = ~new_n14505_ & ~new_n14506_;
  assign new_n14509_ = ~new_n14507_ & new_n14508_;
  assign new_n14510_ = ~new_n14506_ & new_n14507_;
  assign new_n14511_ = new_n4475_ & new_n5074_;
  assign new_n14512_ = ~new_n14505_ & new_n14511_;
  assign new_n14513_ = new_n4219_ & new_n14512_;
  assign new_n14514_ = new_n14510_ & new_n14513_;
  assign new_n14515_ = ~lo0287 & ~new_n4423_;
  assign new_n14516_ = new_n14514_ & new_n14515_;
  assign new_n14517_ = new_n4422_ & new_n14516_;
  assign new_n14518_ = ~new_n14505_ & new_n14506_;
  assign new_n14519_ = ~new_n14507_ & new_n14518_;
  assign new_n14520_ = ~new_n14504_ & ~new_n14509_;
  assign new_n14521_ = ~new_n14517_ & new_n14520_;
  assign li0228 = new_n14519_ | ~new_n14521_;
  assign new_n14523_ = ~new_n3589_ & ~new_n3746_;
  assign new_n14524_ = new_n3740_ & new_n14523_;
  assign new_n14525_ = new_n4024_ & new_n14524_;
  assign new_n14526_ = new_n13448_ & new_n14525_;
  assign new_n14527_ = ~lo0786 & new_n5082_;
  assign new_n14528_ = new_n4422_ & new_n14527_;
  assign new_n14529_ = new_n14515_ & new_n14528_;
  assign new_n14530_ = new_n3612_ & ~new_n14529_;
  assign new_n14531_ = ~new_n3753_ & new_n13457_;
  assign new_n14532_ = new_n3800_ & new_n13453_;
  assign new_n14533_ = ~new_n3763_ & ~new_n4041_;
  assign new_n14534_ = new_n14532_ & new_n14533_;
  assign new_n14535_ = ~new_n3786_ & new_n14534_;
  assign new_n14536_ = ~new_n5562_ & new_n14535_;
  assign new_n14537_ = new_n3917_ & new_n13454_;
  assign new_n14538_ = new_n14536_ & new_n14537_;
  assign new_n14539_ = new_n3941_ & new_n14538_;
  assign new_n14540_ = new_n4117_ & new_n14539_;
  assign new_n14541_ = new_n13463_ & new_n14540_;
  assign new_n14542_ = new_n13482_ & new_n14541_;
  assign new_n14543_ = new_n14526_ & ~new_n14530_;
  assign new_n14544_ = new_n14531_ & new_n14543_;
  assign li0232 = ~new_n14542_ | ~new_n14544_;
  assign new_n14546_ = new_n6057_ & new_n6067_;
  assign new_n14547_ = ~new_n6060_ & new_n14546_;
  assign new_n14548_ = new_n6063_ & new_n14547_;
  assign new_n14549_ = new_n6060_ & ~new_n6063_;
  assign new_n14550_ = new_n14546_ & new_n14549_;
  assign new_n14551_ = new_n6064_ & new_n14546_;
  assign new_n14552_ = ~new_n14548_ & ~new_n14550_;
  assign new_n14553_ = ~new_n14551_ & new_n14552_;
  assign new_n14554_ = ~new_n6060_ & new_n6063_;
  assign new_n14555_ = new_n8536_ & new_n14554_;
  assign new_n14556_ = new_n6060_ & new_n8536_;
  assign new_n14557_ = ~new_n6063_ & new_n14556_;
  assign new_n14558_ = ~new_n14555_ & ~new_n14557_;
  assign new_n14559_ = pi053 & ~new_n14553_;
  assign new_n14560_ = pi054 & ~new_n14558_;
  assign new_n14561_ = ~new_n14559_ & ~new_n14560_;
  assign new_n14562_ = new_n6060_ & new_n6074_;
  assign new_n14563_ = ~new_n6063_ & new_n14562_;
  assign new_n14564_ = pi055 & new_n14563_;
  assign new_n14565_ = pi054 & new_n6075_;
  assign new_n14566_ = ~new_n14564_ & ~new_n14565_;
  assign new_n14567_ = ~new_n6060_ & new_n6074_;
  assign new_n14568_ = new_n6063_ & new_n14567_;
  assign new_n14569_ = new_n6064_ & new_n8536_;
  assign new_n14570_ = pi055 & new_n14568_;
  assign new_n14571_ = pi053 & new_n14569_;
  assign new_n14572_ = ~new_n14570_ & ~new_n14571_;
  assign new_n14573_ = new_n14561_ & new_n14566_;
  assign new_n14574_ = new_n14572_ & new_n14573_;
  assign new_n14575_ = pi065 & new_n14550_;
  assign new_n14576_ = pi066 & new_n14548_;
  assign new_n14577_ = ~new_n14575_ & ~new_n14576_;
  assign new_n14578_ = pi066 & new_n14557_;
  assign new_n14579_ = pi065 & new_n14569_;
  assign new_n14580_ = ~new_n14578_ & ~new_n14579_;
  assign new_n14581_ = pi067 & new_n14563_;
  assign new_n14582_ = pi066 & new_n6075_;
  assign new_n14583_ = ~new_n14581_ & ~new_n14582_;
  assign new_n14584_ = new_n14580_ & new_n14583_;
  assign new_n14585_ = new_n14577_ & new_n14584_;
  assign new_n14586_ = pi067 & new_n14555_;
  assign new_n14587_ = pi064 & new_n14551_;
  assign new_n14588_ = pi068 & new_n14568_;
  assign new_n14589_ = new_n14585_ & ~new_n14586_;
  assign new_n14590_ = ~new_n14587_ & new_n14589_;
  assign new_n14591_ = ~new_n14588_ & new_n14590_;
  assign new_n14592_ = lo0209 & new_n3522_;
  assign new_n14593_ = lo0213 & ~new_n3522_;
  assign new_n14594_ = ~new_n14592_ & ~new_n14593_;
  assign new_n14595_ = ~new_n14574_ & ~new_n14594_;
  assign new_n14596_ = new_n14574_ & ~new_n14591_;
  assign new_n14597_ = ~new_n14595_ & ~new_n14596_;
  assign new_n14598_ = lo0230 & lo0233;
  assign new_n14599_ = ~lo0233 & ~new_n14597_;
  assign li0233 = new_n14598_ | new_n14599_;
  assign new_n14601_ = pi067 & new_n14568_;
  assign new_n14602_ = pi066 & new_n14555_;
  assign new_n14603_ = ~new_n14601_ & ~new_n14602_;
  assign new_n14604_ = pi065 & new_n14548_;
  assign new_n14605_ = new_n14603_ & ~new_n14604_;
  assign new_n14606_ = pi065 & new_n14551_;
  assign new_n14607_ = new_n14584_ & new_n14605_;
  assign new_n14608_ = ~new_n14606_ & new_n14607_;
  assign new_n14609_ = ~new_n14575_ & new_n14608_;
  assign new_n14610_ = pi063 & ~new_n14553_;
  assign new_n14611_ = pi064 & ~new_n14558_;
  assign new_n14612_ = ~new_n14610_ & ~new_n14611_;
  assign new_n14613_ = pi065 & new_n14563_;
  assign new_n14614_ = pi064 & new_n6075_;
  assign new_n14615_ = ~new_n14613_ & ~new_n14614_;
  assign new_n14616_ = pi065 & new_n14568_;
  assign new_n14617_ = pi063 & new_n14569_;
  assign new_n14618_ = ~new_n14616_ & ~new_n14617_;
  assign new_n14619_ = new_n14612_ & new_n14615_;
  assign new_n14620_ = new_n14618_ & new_n14619_;
  assign new_n14621_ = ~new_n14594_ & ~new_n14609_;
  assign new_n14622_ = new_n14609_ & ~new_n14620_;
  assign new_n14623_ = ~new_n14621_ & ~new_n14622_;
  assign new_n14624_ = lo0230 & lo0234;
  assign new_n14625_ = ~lo0234 & ~new_n14623_;
  assign li0234 = new_n14624_ | new_n14625_;
  assign new_n14627_ = pi067 & new_n6075_;
  assign new_n14628_ = ~new_n14576_ & ~new_n14627_;
  assign new_n14629_ = ~new_n14588_ & new_n14628_;
  assign new_n14630_ = ~new_n14586_ & new_n14629_;
  assign new_n14631_ = pi068 & new_n14563_;
  assign new_n14632_ = pi066 & new_n14569_;
  assign new_n14633_ = ~new_n14631_ & ~new_n14632_;
  assign new_n14634_ = pi067 & new_n14557_;
  assign new_n14635_ = pi066 & new_n14550_;
  assign new_n14636_ = ~new_n14634_ & ~new_n14635_;
  assign new_n14637_ = new_n14630_ & new_n14633_;
  assign new_n14638_ = new_n14636_ & new_n14637_;
  assign new_n14639_ = pi066 & new_n14563_;
  assign new_n14640_ = pi065 & new_n6075_;
  assign new_n14641_ = ~new_n14639_ & ~new_n14640_;
  assign new_n14642_ = pi065 & ~new_n14558_;
  assign new_n14643_ = pi064 & ~new_n14552_;
  assign new_n14644_ = ~new_n14642_ & ~new_n14643_;
  assign new_n14645_ = pi066 & new_n14568_;
  assign new_n14646_ = pi064 & new_n14569_;
  assign new_n14647_ = ~new_n14645_ & ~new_n14646_;
  assign new_n14648_ = new_n14641_ & new_n14644_;
  assign new_n14649_ = new_n14647_ & new_n14648_;
  assign new_n14650_ = ~new_n14594_ & ~new_n14638_;
  assign new_n14651_ = new_n14638_ & ~new_n14649_;
  assign new_n14652_ = ~new_n14650_ & ~new_n14651_;
  assign new_n14653_ = lo0230 & lo0235;
  assign new_n14654_ = ~lo0235 & ~new_n14652_;
  assign li0235 = new_n14653_ | new_n14654_;
  assign new_n14656_ = pi054 & ~new_n14553_;
  assign new_n14657_ = pi055 & ~new_n14558_;
  assign new_n14658_ = ~new_n14656_ & ~new_n14657_;
  assign new_n14659_ = pi056 & new_n14563_;
  assign new_n14660_ = pi055 & new_n6075_;
  assign new_n14661_ = ~new_n14659_ & ~new_n14660_;
  assign new_n14662_ = pi056 & new_n14568_;
  assign new_n14663_ = pi054 & new_n14569_;
  assign new_n14664_ = ~new_n14662_ & ~new_n14663_;
  assign new_n14665_ = new_n14658_ & new_n14661_;
  assign new_n14666_ = new_n14664_ & new_n14665_;
  assign new_n14667_ = pi069 & new_n14568_;
  assign new_n14668_ = pi068 & new_n14555_;
  assign new_n14669_ = ~new_n14667_ & ~new_n14668_;
  assign new_n14670_ = pi067 & new_n14548_;
  assign new_n14671_ = new_n14669_ & ~new_n14670_;
  assign new_n14672_ = ~new_n14606_ & ~new_n14627_;
  assign new_n14673_ = new_n14633_ & new_n14671_;
  assign new_n14674_ = new_n14636_ & new_n14673_;
  assign new_n14675_ = new_n14672_ & new_n14674_;
  assign new_n14676_ = ~new_n14594_ & ~new_n14666_;
  assign new_n14677_ = new_n14666_ & ~new_n14675_;
  assign new_n14678_ = ~new_n14676_ & ~new_n14677_;
  assign new_n14679_ = lo0230 & lo0237;
  assign new_n14680_ = ~lo0237 & ~new_n14678_;
  assign li0237 = new_n14679_ | new_n14680_;
  assign new_n14682_ = pi062 & ~new_n14553_;
  assign new_n14683_ = pi063 & ~new_n14558_;
  assign new_n14684_ = ~new_n14682_ & ~new_n14683_;
  assign new_n14685_ = pi064 & new_n14563_;
  assign new_n14686_ = pi063 & new_n6075_;
  assign new_n14687_ = ~new_n14685_ & ~new_n14686_;
  assign new_n14688_ = pi064 & new_n14568_;
  assign new_n14689_ = pi062 & new_n14569_;
  assign new_n14690_ = ~new_n14688_ & ~new_n14689_;
  assign new_n14691_ = new_n14684_ & new_n14687_;
  assign new_n14692_ = new_n14690_ & new_n14691_;
  assign new_n14693_ = ~new_n14587_ & new_n14594_;
  assign new_n14694_ = new_n14649_ & new_n14693_;
  assign new_n14695_ = ~new_n14594_ & new_n14692_;
  assign new_n14696_ = ~new_n14694_ & ~new_n14695_;
  assign new_n14697_ = lo0230 & lo0238;
  assign new_n14698_ = ~lo0238 & new_n14696_;
  assign li0238 = new_n14697_ | new_n14698_;
  assign new_n14700_ = ~new_n14594_ & ~new_n14605_;
  assign new_n14701_ = new_n14594_ & ~new_n14671_;
  assign new_n14702_ = ~new_n14700_ & ~new_n14701_;
  assign new_n14703_ = lo0230 & lo0239;
  assign new_n14704_ = ~lo0239 & ~new_n14702_;
  assign li0239 = new_n14703_ | new_n14704_;
  assign new_n14706_ = pi058 & ~new_n14553_;
  assign new_n14707_ = pi059 & ~new_n14558_;
  assign new_n14708_ = ~new_n14706_ & ~new_n14707_;
  assign new_n14709_ = pi060 & new_n14563_;
  assign new_n14710_ = pi059 & new_n6075_;
  assign new_n14711_ = ~new_n14709_ & ~new_n14710_;
  assign new_n14712_ = pi060 & new_n14568_;
  assign new_n14713_ = pi058 & new_n14569_;
  assign new_n14714_ = ~new_n14712_ & ~new_n14713_;
  assign new_n14715_ = new_n14708_ & new_n14711_;
  assign new_n14716_ = new_n14714_ & new_n14715_;
  assign new_n14717_ = pi056 & ~new_n14553_;
  assign new_n14718_ = pi057 & ~new_n14558_;
  assign new_n14719_ = ~new_n14717_ & ~new_n14718_;
  assign new_n14720_ = pi058 & new_n14563_;
  assign new_n14721_ = pi057 & new_n6075_;
  assign new_n14722_ = ~new_n14720_ & ~new_n14721_;
  assign new_n14723_ = pi058 & new_n14568_;
  assign new_n14724_ = pi056 & new_n14569_;
  assign new_n14725_ = ~new_n14723_ & ~new_n14724_;
  assign new_n14726_ = new_n14719_ & new_n14722_;
  assign new_n14727_ = new_n14725_ & new_n14726_;
  assign new_n14728_ = ~new_n14594_ & ~new_n14716_;
  assign new_n14729_ = new_n14716_ & ~new_n14727_;
  assign new_n14730_ = ~new_n14728_ & ~new_n14729_;
  assign new_n14731_ = lo0230 & lo0240;
  assign new_n14732_ = ~lo0240 & ~new_n14730_;
  assign li0240 = new_n14731_ | new_n14732_;
  assign new_n14734_ = pi060 & ~new_n14553_;
  assign new_n14735_ = pi061 & ~new_n14558_;
  assign new_n14736_ = ~new_n14734_ & ~new_n14735_;
  assign new_n14737_ = pi062 & new_n14563_;
  assign new_n14738_ = pi061 & new_n6075_;
  assign new_n14739_ = ~new_n14737_ & ~new_n14738_;
  assign new_n14740_ = pi062 & new_n14568_;
  assign new_n14741_ = pi060 & new_n14569_;
  assign new_n14742_ = ~new_n14740_ & ~new_n14741_;
  assign new_n14743_ = new_n14736_ & new_n14739_;
  assign new_n14744_ = new_n14742_ & new_n14743_;
  assign new_n14745_ = ~new_n14594_ & ~new_n14692_;
  assign new_n14746_ = new_n14692_ & ~new_n14744_;
  assign new_n14747_ = ~new_n14745_ & ~new_n14746_;
  assign new_n14748_ = lo0230 & lo0241;
  assign new_n14749_ = ~lo0241 & ~new_n14747_;
  assign li0241 = new_n14748_ | new_n14749_;
  assign new_n14751_ = pi055 & ~new_n14553_;
  assign new_n14752_ = pi056 & ~new_n14558_;
  assign new_n14753_ = ~new_n14751_ & ~new_n14752_;
  assign new_n14754_ = pi057 & new_n14563_;
  assign new_n14755_ = pi056 & new_n6075_;
  assign new_n14756_ = ~new_n14754_ & ~new_n14755_;
  assign new_n14757_ = pi057 & new_n14568_;
  assign new_n14758_ = pi055 & new_n14569_;
  assign new_n14759_ = ~new_n14757_ & ~new_n14758_;
  assign new_n14760_ = new_n14753_ & new_n14756_;
  assign new_n14761_ = new_n14759_ & new_n14760_;
  assign new_n14762_ = ~new_n14594_ & ~new_n14761_;
  assign new_n14763_ = ~new_n14574_ & new_n14761_;
  assign new_n14764_ = ~new_n14762_ & ~new_n14763_;
  assign new_n14765_ = lo0230 & lo0242;
  assign new_n14766_ = ~lo0242 & ~new_n14764_;
  assign li0242 = new_n14765_ | new_n14766_;
  assign new_n14768_ = lo0314 & ~new_n3568_;
  assign new_n14769_ = ~new_n6074_ & ~new_n8536_;
  assign new_n14770_ = ~lo0081 & ~lo0085;
  assign new_n14771_ = lo0314 & new_n3568_;
  assign new_n14772_ = ~new_n14769_ & new_n14771_;
  assign new_n14773_ = ~new_n14770_ & new_n14772_;
  assign new_n14774_ = ~new_n14768_ & ~new_n14773_;
  assign new_n14775_ = lo0268 & lo0275;
  assign new_n14776_ = lo0276 & lo0802;
  assign new_n14777_ = lo0271 & new_n14776_;
  assign new_n14778_ = lo0273 & new_n14777_;
  assign new_n14779_ = lo0283 & new_n14778_;
  assign new_n14780_ = new_n14775_ & new_n14779_;
  assign new_n14781_ = lo0272 & new_n14780_;
  assign new_n14782_ = lo0253 & lo0254;
  assign new_n14783_ = new_n14781_ & new_n14782_;
  assign new_n14784_ = lo0263 & new_n14783_;
  assign new_n14785_ = lo0267 & new_n14784_;
  assign new_n14786_ = ~lo0243 & ~new_n14785_;
  assign new_n14787_ = lo0243 & new_n14785_;
  assign new_n14788_ = ~new_n14786_ & ~new_n14787_;
  assign new_n14789_ = ~new_n14774_ & new_n14788_;
  assign new_n14790_ = lo0243 & new_n14774_;
  assign new_n14791_ = ~new_n14789_ & ~new_n14790_;
  assign new_n14792_ = ~pi002 & ~lo0230;
  assign new_n14793_ = ~new_n14791_ & new_n14792_;
  assign new_n14794_ = pi066 & new_n6074_;
  assign new_n14795_ = pi068 & new_n14546_;
  assign new_n14796_ = pi067 & new_n8536_;
  assign new_n14797_ = ~new_n14795_ & ~new_n14796_;
  assign new_n14798_ = ~new_n14794_ & new_n14797_;
  assign new_n14799_ = ~new_n14792_ & ~new_n14798_;
  assign li0243 = new_n14793_ | new_n14799_;
  assign new_n14801_ = ~new_n14594_ & ~new_n14727_;
  assign new_n14802_ = ~new_n14666_ & new_n14727_;
  assign new_n14803_ = ~new_n14801_ & ~new_n14802_;
  assign new_n14804_ = lo0230 & lo0244;
  assign new_n14805_ = ~lo0244 & ~new_n14803_;
  assign li0244 = new_n14804_ | new_n14805_;
  assign new_n14807_ = pi057 & ~new_n14553_;
  assign new_n14808_ = pi058 & ~new_n14558_;
  assign new_n14809_ = ~new_n14807_ & ~new_n14808_;
  assign new_n14810_ = pi059 & new_n14563_;
  assign new_n14811_ = pi058 & new_n6075_;
  assign new_n14812_ = ~new_n14810_ & ~new_n14811_;
  assign new_n14813_ = pi059 & new_n14568_;
  assign new_n14814_ = pi057 & new_n14569_;
  assign new_n14815_ = ~new_n14813_ & ~new_n14814_;
  assign new_n14816_ = new_n14809_ & new_n14812_;
  assign new_n14817_ = new_n14815_ & new_n14816_;
  assign new_n14818_ = ~new_n14594_ & ~new_n14817_;
  assign new_n14819_ = ~new_n14761_ & new_n14817_;
  assign new_n14820_ = ~new_n14818_ & ~new_n14819_;
  assign new_n14821_ = lo0230 & lo0245;
  assign new_n14822_ = ~lo0245 & ~new_n14820_;
  assign li0245 = new_n14821_ | new_n14822_;
  assign new_n14824_ = pi059 & ~new_n14553_;
  assign new_n14825_ = pi060 & ~new_n14558_;
  assign new_n14826_ = ~new_n14824_ & ~new_n14825_;
  assign new_n14827_ = pi061 & new_n14563_;
  assign new_n14828_ = pi060 & new_n6075_;
  assign new_n14829_ = ~new_n14827_ & ~new_n14828_;
  assign new_n14830_ = pi061 & new_n14568_;
  assign new_n14831_ = pi059 & new_n14569_;
  assign new_n14832_ = ~new_n14830_ & ~new_n14831_;
  assign new_n14833_ = new_n14826_ & new_n14829_;
  assign new_n14834_ = new_n14832_ & new_n14833_;
  assign new_n14835_ = ~new_n14594_ & ~new_n14834_;
  assign new_n14836_ = ~new_n14817_ & new_n14834_;
  assign new_n14837_ = ~new_n14835_ & ~new_n14836_;
  assign new_n14838_ = lo0230 & lo0246;
  assign new_n14839_ = ~lo0246 & ~new_n14837_;
  assign li0246 = new_n14838_ | new_n14839_;
  assign new_n14841_ = ~new_n14594_ & ~new_n14744_;
  assign new_n14842_ = ~new_n14716_ & new_n14744_;
  assign new_n14843_ = ~new_n14841_ & ~new_n14842_;
  assign new_n14844_ = lo0230 & lo0247;
  assign new_n14845_ = ~lo0247 & ~new_n14843_;
  assign li0247 = new_n14844_ | new_n14845_;
  assign new_n14847_ = pi061 & ~new_n14553_;
  assign new_n14848_ = pi062 & ~new_n14558_;
  assign new_n14849_ = ~new_n14847_ & ~new_n14848_;
  assign new_n14850_ = pi063 & new_n14563_;
  assign new_n14851_ = pi062 & new_n6075_;
  assign new_n14852_ = ~new_n14850_ & ~new_n14851_;
  assign new_n14853_ = pi063 & new_n14568_;
  assign new_n14854_ = pi061 & new_n14569_;
  assign new_n14855_ = ~new_n14853_ & ~new_n14854_;
  assign new_n14856_ = new_n14849_ & new_n14852_;
  assign new_n14857_ = new_n14855_ & new_n14856_;
  assign new_n14858_ = ~new_n14594_ & ~new_n14857_;
  assign new_n14859_ = ~new_n14834_ & new_n14857_;
  assign new_n14860_ = ~new_n14858_ & ~new_n14859_;
  assign new_n14861_ = lo0230 & lo0248;
  assign new_n14862_ = ~lo0248 & ~new_n14860_;
  assign li0248 = new_n14861_ | new_n14862_;
  assign new_n14864_ = ~new_n14594_ & ~new_n14620_;
  assign new_n14865_ = new_n14620_ & ~new_n14857_;
  assign new_n14866_ = ~new_n14864_ & ~new_n14865_;
  assign new_n14867_ = lo0230 & lo0249;
  assign new_n14868_ = ~lo0249 & ~new_n14866_;
  assign li0249 = new_n14867_ | new_n14868_;
  assign new_n14870_ = ~new_n3705_ & ~new_n4050_;
  assign new_n14871_ = ~lo0250 & ~new_n13463_;
  assign new_n14872_ = ~lo0250 & new_n13463_;
  assign new_n14873_ = new_n14870_ & ~new_n14872_;
  assign new_n14874_ = ~new_n14871_ & new_n14872_;
  assign new_n14875_ = ~new_n14873_ & ~new_n14874_;
  assign new_n14876_ = ~new_n14870_ & new_n14871_;
  assign li0250 = new_n14875_ | new_n14876_;
  assign new_n14878_ = ~lo0199 & lo0200;
  assign new_n14879_ = lo0476 & new_n14878_;
  assign new_n14880_ = lo1033 & ~new_n14879_;
  assign new_n14881_ = lo0251 & ~lo1033;
  assign new_n14882_ = ~new_n14880_ & ~new_n14881_;
  assign new_n14883_ = ~lo0199 & ~lo0200;
  assign new_n14884_ = lo0897 & new_n14883_;
  assign new_n14885_ = lo1047 & ~new_n14884_;
  assign new_n14886_ = ~lo1047 & ~new_n14882_;
  assign li0251 = new_n14885_ | new_n14886_;
  assign new_n14888_ = pi004 & ~new_n5051_;
  assign new_n14889_ = pi003 & ~new_n14888_;
  assign new_n14890_ = lo0252 & new_n14889_;
  assign new_n14891_ = new_n4475_ & new_n5070_;
  assign li0252 = new_n14890_ | new_n14891_;
  assign new_n14893_ = ~lo0253 & ~new_n14781_;
  assign new_n14894_ = lo0253 & new_n14781_;
  assign new_n14895_ = ~new_n14893_ & ~new_n14894_;
  assign new_n14896_ = ~new_n14774_ & new_n14895_;
  assign new_n14897_ = lo0253 & new_n14774_;
  assign new_n14898_ = ~new_n14896_ & ~new_n14897_;
  assign new_n14899_ = new_n14792_ & ~new_n14898_;
  assign new_n14900_ = pi062 & new_n6074_;
  assign new_n14901_ = pi064 & new_n14546_;
  assign new_n14902_ = pi063 & new_n8536_;
  assign new_n14903_ = ~new_n14901_ & ~new_n14902_;
  assign new_n14904_ = ~new_n14900_ & new_n14903_;
  assign new_n14905_ = ~new_n14792_ & ~new_n14904_;
  assign li0253 = new_n14899_ | new_n14905_;
  assign new_n14907_ = lo0272 & lo0275;
  assign new_n14908_ = lo0253 & lo0268;
  assign new_n14909_ = new_n14907_ & new_n14908_;
  assign new_n14910_ = new_n14779_ & new_n14909_;
  assign new_n14911_ = ~lo0254 & ~new_n14910_;
  assign new_n14912_ = lo0254 & new_n14910_;
  assign new_n14913_ = ~new_n14911_ & ~new_n14912_;
  assign new_n14914_ = ~new_n14774_ & new_n14913_;
  assign new_n14915_ = lo0254 & new_n14774_;
  assign new_n14916_ = ~new_n14914_ & ~new_n14915_;
  assign new_n14917_ = new_n14792_ & ~new_n14916_;
  assign new_n14918_ = pi063 & new_n6074_;
  assign new_n14919_ = pi065 & new_n14546_;
  assign new_n14920_ = pi064 & new_n8536_;
  assign new_n14921_ = ~new_n14919_ & ~new_n14920_;
  assign new_n14922_ = ~new_n14918_ & new_n14921_;
  assign new_n14923_ = ~new_n14792_ & ~new_n14922_;
  assign li0254 = new_n14917_ | new_n14923_;
  assign new_n14925_ = lo1030 & ~new_n14879_;
  assign new_n14926_ = lo0255 & ~lo1030;
  assign new_n14927_ = ~new_n14925_ & ~new_n14926_;
  assign new_n14928_ = lo1043 & ~new_n14884_;
  assign new_n14929_ = ~lo1043 & ~new_n14927_;
  assign li0255 = new_n14928_ | new_n14929_;
  assign new_n14931_ = lo1064 & ~new_n14879_;
  assign new_n14932_ = lo0256 & ~lo1064;
  assign new_n14933_ = ~new_n14931_ & ~new_n14932_;
  assign new_n14934_ = lo1042 & ~new_n14884_;
  assign new_n14935_ = ~lo1042 & ~new_n14933_;
  assign li0256 = new_n14934_ | new_n14935_;
  assign new_n14937_ = lo1059 & ~new_n14879_;
  assign new_n14938_ = lo0257 & ~lo1059;
  assign new_n14939_ = ~new_n14937_ & ~new_n14938_;
  assign new_n14940_ = lo1078 & ~new_n14884_;
  assign new_n14941_ = ~lo1078 & ~new_n14939_;
  assign li0257 = new_n14940_ | new_n14941_;
  assign new_n14943_ = lo1056 & ~new_n14879_;
  assign new_n14944_ = lo0258 & ~lo1056;
  assign new_n14945_ = ~new_n14943_ & ~new_n14944_;
  assign new_n14946_ = lo1066 & ~new_n14884_;
  assign new_n14947_ = ~lo1066 & ~new_n14945_;
  assign li0258 = new_n14946_ | new_n14947_;
  assign new_n14949_ = lo1063 & ~new_n14879_;
  assign new_n14950_ = lo0259 & ~lo1063;
  assign new_n14951_ = ~new_n14949_ & ~new_n14950_;
  assign new_n14952_ = lo1053 & ~new_n14884_;
  assign new_n14953_ = ~lo1053 & ~new_n14951_;
  assign li0259 = new_n14952_ | new_n14953_;
  assign new_n14955_ = lo1061 & ~new_n14879_;
  assign new_n14956_ = lo0260 & ~lo1061;
  assign new_n14957_ = ~new_n14955_ & ~new_n14956_;
  assign new_n14958_ = lo1038 & ~new_n14884_;
  assign new_n14959_ = ~lo1038 & ~new_n14957_;
  assign li0260 = new_n14958_ | new_n14959_;
  assign new_n14961_ = lo1034 & ~new_n14879_;
  assign new_n14962_ = lo0261 & ~lo1034;
  assign new_n14963_ = ~new_n14961_ & ~new_n14962_;
  assign new_n14964_ = lo1031 & ~new_n14884_;
  assign new_n14965_ = ~lo1031 & ~new_n14963_;
  assign li0261 = new_n14964_ | new_n14965_;
  assign new_n14967_ = ~new_n14557_ & ~new_n14563_;
  assign new_n14968_ = ~new_n6075_ & new_n14967_;
  assign new_n14969_ = ~new_n14555_ & ~new_n14568_;
  assign new_n14970_ = pi053 & ~new_n14968_;
  assign new_n14971_ = pi053 & ~new_n14969_;
  assign new_n14972_ = ~new_n14970_ & ~new_n14971_;
  assign new_n14973_ = lo0123 & ~lo0228;
  assign new_n14974_ = pi004 & ~lo0123;
  assign new_n14975_ = ~new_n14973_ & ~new_n14974_;
  assign new_n14976_ = lo0262 & new_n14975_;
  assign new_n14977_ = ~new_n14972_ & ~new_n14975_;
  assign li0262 = new_n14976_ | new_n14977_;
  assign new_n14979_ = new_n14779_ & new_n14907_;
  assign new_n14980_ = new_n14908_ & new_n14979_;
  assign new_n14981_ = lo0267 & new_n14980_;
  assign new_n14982_ = lo0254 & new_n14981_;
  assign new_n14983_ = ~lo0263 & ~new_n14982_;
  assign new_n14984_ = lo0263 & new_n14982_;
  assign new_n14985_ = ~new_n14983_ & ~new_n14984_;
  assign new_n14986_ = ~new_n14774_ & new_n14985_;
  assign new_n14987_ = lo0263 & new_n14774_;
  assign new_n14988_ = ~new_n14986_ & ~new_n14987_;
  assign new_n14989_ = new_n14792_ & ~new_n14988_;
  assign new_n14990_ = pi065 & new_n6074_;
  assign new_n14991_ = pi067 & new_n14546_;
  assign new_n14992_ = pi066 & new_n8536_;
  assign new_n14993_ = ~new_n14991_ & ~new_n14992_;
  assign new_n14994_ = ~new_n14990_ & new_n14993_;
  assign new_n14995_ = ~new_n14792_ & ~new_n14994_;
  assign li0263 = new_n14989_ | new_n14995_;
  assign new_n14997_ = lo0796 & new_n14774_;
  assign new_n14998_ = lo0264 & ~lo0796;
  assign new_n14999_ = ~new_n14997_ & ~new_n14998_;
  assign new_n15000_ = pi052 & new_n6074_;
  assign new_n15001_ = pi054 & new_n14546_;
  assign new_n15002_ = pi053 & new_n8536_;
  assign new_n15003_ = ~new_n15001_ & ~new_n15002_;
  assign new_n15004_ = ~new_n15000_ & new_n15003_;
  assign new_n15005_ = ~new_n14792_ & ~new_n15004_;
  assign new_n15006_ = new_n14792_ & ~new_n14999_;
  assign li0264 = new_n15005_ | new_n15006_;
  assign new_n15008_ = lo0819 & new_n14774_;
  assign new_n15009_ = lo0265 & ~lo0819;
  assign new_n15010_ = ~new_n15008_ & ~new_n15009_;
  assign new_n15011_ = pi053 & new_n6074_;
  assign new_n15012_ = pi055 & new_n14546_;
  assign new_n15013_ = pi054 & new_n8536_;
  assign new_n15014_ = ~new_n15012_ & ~new_n15013_;
  assign new_n15015_ = ~new_n15011_ & new_n15014_;
  assign new_n15016_ = ~new_n14792_ & ~new_n15015_;
  assign new_n15017_ = new_n14792_ & ~new_n15010_;
  assign li0265 = new_n15016_ | new_n15017_;
  assign new_n15019_ = lo0948 & new_n14774_;
  assign new_n15020_ = lo0266 & ~lo0948;
  assign new_n15021_ = ~new_n15019_ & ~new_n15020_;
  assign new_n15022_ = pi045 & new_n6074_;
  assign new_n15023_ = pi047 & new_n14546_;
  assign new_n15024_ = pi046 & new_n8536_;
  assign new_n15025_ = ~new_n15023_ & ~new_n15024_;
  assign new_n15026_ = ~new_n15022_ & new_n15025_;
  assign new_n15027_ = ~new_n14792_ & ~new_n15026_;
  assign new_n15028_ = new_n14792_ & ~new_n15021_;
  assign li0266 = new_n15027_ | new_n15028_;
  assign new_n15030_ = pi066 & new_n14546_;
  assign new_n15031_ = pi065 & new_n8536_;
  assign new_n15032_ = ~new_n15030_ & ~new_n15031_;
  assign new_n15033_ = pi064 & new_n6074_;
  assign new_n15034_ = new_n15032_ & ~new_n15033_;
  assign new_n15035_ = lo0271 & lo0273;
  assign new_n15036_ = lo0272 & new_n15035_;
  assign new_n15037_ = lo0283 & new_n15036_;
  assign new_n15038_ = new_n14776_ & new_n15037_;
  assign new_n15039_ = new_n14775_ & new_n15038_;
  assign new_n15040_ = new_n14782_ & new_n15039_;
  assign new_n15041_ = ~lo0267 & ~new_n15040_;
  assign new_n15042_ = lo0267 & new_n15040_;
  assign new_n15043_ = ~new_n15041_ & ~new_n15042_;
  assign new_n15044_ = ~new_n14774_ & new_n15043_;
  assign new_n15045_ = lo0267 & new_n14774_;
  assign new_n15046_ = ~new_n15044_ & ~new_n15045_;
  assign new_n15047_ = ~new_n14792_ & ~new_n15034_;
  assign new_n15048_ = new_n14792_ & ~new_n15046_;
  assign li0267 = new_n15047_ | new_n15048_;
  assign new_n15050_ = ~lo0268 & new_n14979_;
  assign new_n15051_ = lo0268 & ~new_n14979_;
  assign new_n15052_ = ~new_n15050_ & ~new_n15051_;
  assign new_n15053_ = new_n14774_ & ~new_n15052_;
  assign new_n15054_ = lo0268 & new_n15052_;
  assign new_n15055_ = ~new_n15053_ & ~new_n15054_;
  assign new_n15056_ = pi061 & new_n6074_;
  assign new_n15057_ = pi063 & new_n14546_;
  assign new_n15058_ = pi062 & new_n8536_;
  assign new_n15059_ = ~new_n15057_ & ~new_n15058_;
  assign new_n15060_ = ~new_n15056_ & new_n15059_;
  assign new_n15061_ = ~new_n14792_ & ~new_n15060_;
  assign new_n15062_ = new_n14792_ & ~new_n15055_;
  assign li0268 = new_n15061_ | new_n15062_;
  assign new_n15064_ = lo0817 & new_n14774_;
  assign new_n15065_ = lo0269 & ~lo0817;
  assign new_n15066_ = ~new_n15064_ & ~new_n15065_;
  assign new_n15067_ = pi047 & new_n6074_;
  assign new_n15068_ = pi049 & new_n14546_;
  assign new_n15069_ = pi048 & new_n8536_;
  assign new_n15070_ = ~new_n15068_ & ~new_n15069_;
  assign new_n15071_ = ~new_n15067_ & new_n15070_;
  assign new_n15072_ = ~new_n14792_ & ~new_n15071_;
  assign new_n15073_ = new_n14792_ & ~new_n15066_;
  assign li0269 = new_n15072_ | new_n15073_;
  assign new_n15075_ = lo0805 & new_n14774_;
  assign new_n15076_ = lo0270 & ~lo0805;
  assign new_n15077_ = ~new_n15075_ & ~new_n15076_;
  assign new_n15078_ = pi050 & new_n6074_;
  assign new_n15079_ = pi052 & new_n14546_;
  assign new_n15080_ = pi051 & new_n8536_;
  assign new_n15081_ = ~new_n15079_ & ~new_n15080_;
  assign new_n15082_ = ~new_n15078_ & new_n15081_;
  assign new_n15083_ = ~new_n14792_ & ~new_n15082_;
  assign new_n15084_ = new_n14792_ & ~new_n15077_;
  assign li0270 = new_n15083_ | new_n15084_;
  assign new_n15086_ = ~lo0271 & new_n14776_;
  assign new_n15087_ = lo0271 & ~new_n14776_;
  assign new_n15088_ = ~new_n15086_ & ~new_n15087_;
  assign new_n15089_ = new_n14774_ & ~new_n15088_;
  assign new_n15090_ = lo0271 & new_n15088_;
  assign new_n15091_ = ~new_n15089_ & ~new_n15090_;
  assign new_n15092_ = pi056 & new_n6074_;
  assign new_n15093_ = pi058 & new_n14546_;
  assign new_n15094_ = pi057 & new_n8536_;
  assign new_n15095_ = ~new_n15093_ & ~new_n15094_;
  assign new_n15096_ = ~new_n15092_ & new_n15095_;
  assign new_n15097_ = ~new_n14792_ & ~new_n15096_;
  assign new_n15098_ = new_n14792_ & ~new_n15091_;
  assign li0271 = new_n15097_ | new_n15098_;
  assign new_n15100_ = ~lo0272 & new_n14779_;
  assign new_n15101_ = lo0272 & ~new_n14779_;
  assign new_n15102_ = ~new_n15100_ & ~new_n15101_;
  assign new_n15103_ = new_n14774_ & ~new_n15102_;
  assign new_n15104_ = lo0272 & new_n15102_;
  assign new_n15105_ = ~new_n15103_ & ~new_n15104_;
  assign new_n15106_ = pi059 & new_n6074_;
  assign new_n15107_ = pi061 & new_n14546_;
  assign new_n15108_ = pi060 & new_n8536_;
  assign new_n15109_ = ~new_n15107_ & ~new_n15108_;
  assign new_n15110_ = ~new_n15106_ & new_n15109_;
  assign new_n15111_ = ~new_n14792_ & ~new_n15110_;
  assign new_n15112_ = new_n14792_ & ~new_n15105_;
  assign li0272 = new_n15111_ | new_n15112_;
  assign new_n15114_ = ~lo0273 & new_n14777_;
  assign new_n15115_ = lo0273 & ~new_n14777_;
  assign new_n15116_ = ~new_n15114_ & ~new_n15115_;
  assign new_n15117_ = new_n14774_ & ~new_n15116_;
  assign new_n15118_ = lo0273 & new_n15116_;
  assign new_n15119_ = ~new_n15117_ & ~new_n15118_;
  assign new_n15120_ = pi057 & new_n6074_;
  assign new_n15121_ = pi059 & new_n14546_;
  assign new_n15122_ = pi058 & new_n8536_;
  assign new_n15123_ = ~new_n15121_ & ~new_n15122_;
  assign new_n15124_ = ~new_n15120_ & new_n15123_;
  assign new_n15125_ = ~new_n14792_ & ~new_n15124_;
  assign new_n15126_ = new_n14792_ & ~new_n15119_;
  assign li0273 = new_n15125_ | new_n15126_;
  assign new_n15128_ = lo0659 & new_n14774_;
  assign new_n15129_ = lo0274 & ~lo0659;
  assign new_n15130_ = ~new_n15128_ & ~new_n15129_;
  assign new_n15131_ = pi054 & new_n6074_;
  assign new_n15132_ = pi056 & new_n14546_;
  assign new_n15133_ = pi055 & new_n8536_;
  assign new_n15134_ = ~new_n15132_ & ~new_n15133_;
  assign new_n15135_ = ~new_n15131_ & new_n15134_;
  assign new_n15136_ = ~new_n14792_ & ~new_n15135_;
  assign new_n15137_ = new_n14792_ & ~new_n15130_;
  assign li0274 = new_n15136_ | new_n15137_;
  assign new_n15139_ = ~lo0275 & new_n15038_;
  assign new_n15140_ = lo0275 & ~new_n15038_;
  assign new_n15141_ = ~new_n15139_ & ~new_n15140_;
  assign new_n15142_ = new_n14774_ & ~new_n15141_;
  assign new_n15143_ = lo0275 & new_n15141_;
  assign new_n15144_ = ~new_n15142_ & ~new_n15143_;
  assign new_n15145_ = pi060 & new_n6074_;
  assign new_n15146_ = pi062 & new_n14546_;
  assign new_n15147_ = pi061 & new_n8536_;
  assign new_n15148_ = ~new_n15146_ & ~new_n15147_;
  assign new_n15149_ = ~new_n15145_ & new_n15148_;
  assign new_n15150_ = ~new_n14792_ & ~new_n15149_;
  assign new_n15151_ = new_n14792_ & ~new_n15144_;
  assign li0275 = new_n15150_ | new_n15151_;
  assign new_n15153_ = lo0276 & ~lo0802;
  assign new_n15154_ = ~lo0276 & lo0802;
  assign new_n15155_ = ~new_n15153_ & ~new_n15154_;
  assign new_n15156_ = new_n14774_ & ~new_n15155_;
  assign new_n15157_ = lo0276 & new_n15155_;
  assign new_n15158_ = ~new_n15156_ & ~new_n15157_;
  assign new_n15159_ = pi055 & new_n6074_;
  assign new_n15160_ = pi057 & new_n14546_;
  assign new_n15161_ = pi056 & new_n8536_;
  assign new_n15162_ = ~new_n15160_ & ~new_n15161_;
  assign new_n15163_ = ~new_n15159_ & new_n15162_;
  assign new_n15164_ = ~new_n14792_ & ~new_n15163_;
  assign new_n15165_ = new_n14792_ & ~new_n15158_;
  assign li0276 = new_n15164_ | new_n15165_;
  assign new_n15167_ = lo0820 & new_n14774_;
  assign new_n15168_ = lo0277 & ~lo0820;
  assign new_n15169_ = ~new_n15167_ & ~new_n15168_;
  assign new_n15170_ = pi051 & new_n6074_;
  assign new_n15171_ = pi053 & new_n14546_;
  assign new_n15172_ = pi052 & new_n8536_;
  assign new_n15173_ = ~new_n15171_ & ~new_n15172_;
  assign new_n15174_ = ~new_n15170_ & new_n15173_;
  assign new_n15175_ = ~new_n14792_ & ~new_n15174_;
  assign new_n15176_ = new_n14792_ & ~new_n15169_;
  assign li0277 = new_n15175_ | new_n15176_;
  assign new_n15178_ = lo0976 & new_n14774_;
  assign new_n15179_ = lo0278 & ~lo0976;
  assign new_n15180_ = ~new_n15178_ & ~new_n15179_;
  assign new_n15181_ = pi045 & new_n14546_;
  assign new_n15182_ = pi043 & new_n6074_;
  assign new_n15183_ = pi044 & new_n8536_;
  assign new_n15184_ = ~new_n15182_ & ~new_n15183_;
  assign new_n15185_ = ~new_n15181_ & new_n15184_;
  assign new_n15186_ = ~new_n14792_ & ~new_n15185_;
  assign new_n15187_ = new_n14792_ & ~new_n15180_;
  assign li0278 = new_n15186_ | new_n15187_;
  assign new_n15189_ = lo0958 & new_n14774_;
  assign new_n15190_ = lo0279 & ~lo0958;
  assign new_n15191_ = ~new_n15189_ & ~new_n15190_;
  assign new_n15192_ = pi045 & new_n8536_;
  assign new_n15193_ = pi044 & new_n6074_;
  assign new_n15194_ = pi046 & new_n14546_;
  assign new_n15195_ = ~new_n15193_ & ~new_n15194_;
  assign new_n15196_ = ~new_n15192_ & new_n15195_;
  assign new_n15197_ = ~new_n14792_ & ~new_n15196_;
  assign new_n15198_ = new_n14792_ & ~new_n15191_;
  assign li0279 = new_n15197_ | new_n15198_;
  assign new_n15200_ = lo0914 & new_n14774_;
  assign new_n15201_ = lo0280 & ~lo0914;
  assign new_n15202_ = ~new_n15200_ & ~new_n15201_;
  assign new_n15203_ = pi046 & new_n6074_;
  assign new_n15204_ = pi048 & new_n14546_;
  assign new_n15205_ = pi047 & new_n8536_;
  assign new_n15206_ = ~new_n15204_ & ~new_n15205_;
  assign new_n15207_ = ~new_n15203_ & new_n15206_;
  assign new_n15208_ = ~new_n14792_ & ~new_n15207_;
  assign new_n15209_ = new_n14792_ & ~new_n15202_;
  assign li0280 = new_n15208_ | new_n15209_;
  assign new_n15211_ = lo0830 & new_n14774_;
  assign new_n15212_ = lo0281 & ~lo0830;
  assign new_n15213_ = ~new_n15211_ & ~new_n15212_;
  assign new_n15214_ = pi048 & new_n6074_;
  assign new_n15215_ = pi050 & new_n14546_;
  assign new_n15216_ = pi049 & new_n8536_;
  assign new_n15217_ = ~new_n15215_ & ~new_n15216_;
  assign new_n15218_ = ~new_n15214_ & new_n15217_;
  assign new_n15219_ = ~new_n14792_ & ~new_n15218_;
  assign new_n15220_ = new_n14792_ & ~new_n15213_;
  assign li0281 = new_n15219_ | new_n15220_;
  assign new_n15222_ = lo0836 & new_n14774_;
  assign new_n15223_ = lo0282 & ~lo0836;
  assign new_n15224_ = ~new_n15222_ & ~new_n15223_;
  assign new_n15225_ = pi049 & new_n6074_;
  assign new_n15226_ = pi051 & new_n14546_;
  assign new_n15227_ = pi050 & new_n8536_;
  assign new_n15228_ = ~new_n15226_ & ~new_n15227_;
  assign new_n15229_ = ~new_n15225_ & new_n15228_;
  assign new_n15230_ = ~new_n14792_ & ~new_n15229_;
  assign new_n15231_ = new_n14792_ & ~new_n15224_;
  assign li0282 = new_n15230_ | new_n15231_;
  assign new_n15233_ = ~lo0283 & new_n14778_;
  assign new_n15234_ = lo0283 & ~new_n14778_;
  assign new_n15235_ = ~new_n15233_ & ~new_n15234_;
  assign new_n15236_ = new_n14774_ & ~new_n15235_;
  assign new_n15237_ = lo0283 & new_n15235_;
  assign new_n15238_ = ~new_n15236_ & ~new_n15237_;
  assign new_n15239_ = pi058 & new_n6074_;
  assign new_n15240_ = pi060 & new_n14546_;
  assign new_n15241_ = pi059 & new_n8536_;
  assign new_n15242_ = ~new_n15240_ & ~new_n15241_;
  assign new_n15243_ = ~new_n15239_ & new_n15242_;
  assign new_n15244_ = ~new_n14792_ & ~new_n15243_;
  assign new_n15245_ = new_n14792_ & ~new_n15238_;
  assign li0283 = new_n15244_ | new_n15245_;
  assign new_n15247_ = pi054 & ~new_n14975_;
  assign new_n15248_ = ~new_n14563_ & ~new_n14568_;
  assign new_n15249_ = new_n15247_ & ~new_n15248_;
  assign new_n15250_ = lo0284 & new_n14975_;
  assign li0284 = new_n15249_ | new_n15250_;
  assign new_n15252_ = lo0286 & lo0288;
  assign new_n15253_ = lo0289 & new_n15252_;
  assign new_n15254_ = ~lo0285 & ~new_n15253_;
  assign new_n15255_ = lo0285 & new_n15253_;
  assign new_n15256_ = ~new_n15254_ & ~new_n15255_;
  assign new_n15257_ = lo0285 & ~new_n4668_;
  assign new_n15258_ = ~new_n4669_ & ~new_n15257_;
  assign new_n15259_ = new_n4672_ & ~li0480;
  assign new_n15260_ = ~lo0285 & new_n15259_;
  assign new_n15261_ = lo0285 & new_n15258_;
  assign new_n15262_ = ~new_n15260_ & ~new_n15261_;
  assign new_n15263_ = ~new_n4672_ & li0480;
  assign new_n15264_ = ~new_n15256_ & ~new_n15263_;
  assign new_n15265_ = new_n15256_ & ~new_n15262_;
  assign new_n15266_ = ~new_n15264_ & ~new_n15265_;
  assign li0285 = ~lo0793 & new_n15266_;
  assign new_n15268_ = ~new_n4667_ & ~new_n15252_;
  assign new_n15269_ = lo0286 & new_n15259_;
  assign new_n15270_ = ~lo0286 & ~new_n15268_;
  assign new_n15271_ = ~new_n15269_ & ~new_n15270_;
  assign new_n15272_ = ~lo0286 & lo0288;
  assign new_n15273_ = lo0286 & ~lo0288;
  assign new_n15274_ = ~new_n15272_ & ~new_n15273_;
  assign new_n15275_ = ~new_n15263_ & ~new_n15271_;
  assign new_n15276_ = new_n15263_ & ~new_n15274_;
  assign new_n15277_ = ~new_n15275_ & ~new_n15276_;
  assign li0286 = ~lo0793 & ~new_n15277_;
  assign new_n15279_ = ~lo0287 & ~lo0457;
  assign li0287 = ~lo0332 & ~new_n15279_;
  assign new_n15281_ = ~lo0288 & new_n15259_;
  assign new_n15282_ = lo0288 & ~new_n15259_;
  assign new_n15283_ = ~new_n15281_ & ~new_n15282_;
  assign new_n15284_ = ~lo0288 & new_n15263_;
  assign new_n15285_ = ~new_n15263_ & ~new_n15283_;
  assign new_n15286_ = ~new_n15284_ & ~new_n15285_;
  assign li0288 = ~lo0793 & ~new_n15286_;
  assign new_n15288_ = ~lo0289 & ~new_n15252_;
  assign new_n15289_ = ~new_n15253_ & ~new_n15288_;
  assign new_n15290_ = lo0289 & ~new_n4667_;
  assign new_n15291_ = ~new_n4668_ & ~new_n15290_;
  assign new_n15292_ = ~lo0289 & new_n15259_;
  assign new_n15293_ = lo0289 & new_n15291_;
  assign new_n15294_ = ~new_n15292_ & ~new_n15293_;
  assign new_n15295_ = ~new_n15263_ & ~new_n15289_;
  assign new_n15296_ = new_n15289_ & ~new_n15294_;
  assign new_n15297_ = ~new_n15295_ & ~new_n15296_;
  assign li0289 = ~lo0793 & new_n15297_;
  assign new_n15299_ = ~lo0476 & lo1042;
  assign new_n15300_ = lo0290 & ~lo1042;
  assign li0290 = new_n15299_ | new_n15300_;
  assign new_n15302_ = ~lo0476 & lo1043;
  assign new_n15303_ = lo0291 & ~lo1043;
  assign li0291 = new_n15302_ | new_n15303_;
  assign new_n15305_ = ~lo0476 & lo1078;
  assign new_n15306_ = lo0292 & ~lo1078;
  assign li0292 = new_n15305_ | new_n15306_;
  assign new_n15308_ = ~lo0476 & lo1053;
  assign new_n15309_ = lo0293 & ~lo1053;
  assign li0293 = new_n15308_ | new_n15309_;
  assign new_n15311_ = ~lo0476 & lo1066;
  assign new_n15312_ = lo0294 & ~lo1066;
  assign li0294 = new_n15311_ | new_n15312_;
  assign new_n15314_ = ~lo0476 & lo1047;
  assign new_n15315_ = lo0295 & ~lo1047;
  assign li0295 = new_n15314_ | new_n15315_;
  assign new_n15317_ = ~lo0476 & lo1031;
  assign new_n15318_ = lo0296 & ~lo1031;
  assign li0296 = new_n15317_ | new_n15318_;
  assign new_n15320_ = ~lo0476 & lo1038;
  assign new_n15321_ = lo0297 & ~lo1038;
  assign li0297 = new_n15320_ | new_n15321_;
  assign new_n15323_ = ~lo0478 & lo1038;
  assign new_n15324_ = lo0298 & ~lo1038;
  assign li0298 = new_n15323_ | new_n15324_;
  assign new_n15326_ = lo0039 & new_n6962_;
  assign new_n15327_ = new_n14260_ & new_n14266_;
  assign new_n15328_ = new_n3842_ & new_n13346_;
  assign new_n15329_ = ~lo0087 & new_n4171_;
  assign new_n15330_ = new_n14228_ & new_n15329_;
  assign new_n15331_ = new_n4176_ & new_n15330_;
  assign new_n15332_ = new_n14225_ & new_n15331_;
  assign new_n15333_ = new_n15328_ & new_n15332_;
  assign new_n15334_ = new_n4178_ & new_n15333_;
  assign new_n15335_ = ~lo0066 & new_n15334_;
  assign new_n15336_ = ~li0893 & new_n15335_;
  assign new_n15337_ = new_n14224_ & new_n15336_;
  assign new_n15338_ = new_n4154_ & new_n13359_;
  assign new_n15339_ = new_n15337_ & new_n15338_;
  assign new_n15340_ = new_n13344_ & new_n15339_;
  assign new_n15341_ = new_n4153_ & new_n15340_;
  assign new_n15342_ = ~new_n3964_ & ~new_n4130_;
  assign new_n15343_ = new_n15341_ & ~new_n15342_;
  assign new_n15344_ = new_n14255_ & new_n15341_;
  assign new_n15345_ = ~lo0053 & new_n15343_;
  assign new_n15346_ = ~new_n15344_ & ~new_n15345_;
  assign new_n15347_ = new_n15327_ & ~new_n15346_;
  assign new_n15348_ = new_n3535_ & new_n15347_;
  assign new_n15349_ = new_n14262_ & new_n15348_;
  assign new_n15350_ = ~lo0039 & new_n15349_;
  assign new_n15351_ = new_n14268_ & new_n15350_;
  assign li0299 = new_n15326_ | new_n15351_;
  assign new_n15353_ = ~lo0300 & ~lo0312;
  assign new_n15354_ = lo0300 & lo0312;
  assign new_n15355_ = ~new_n15353_ & ~new_n15354_;
  assign new_n15356_ = new_n8092_ & ~new_n15355_;
  assign new_n15357_ = lo0300 & ~new_n8092_;
  assign new_n15358_ = ~new_n15356_ & ~new_n15357_;
  assign li0300 = lo0055 | ~new_n15358_;
  assign new_n15360_ = ~lo0301 & new_n15353_;
  assign new_n15361_ = lo0301 & ~new_n15353_;
  assign new_n15362_ = ~new_n15360_ & ~new_n15361_;
  assign new_n15363_ = new_n8092_ & ~new_n15362_;
  assign new_n15364_ = lo0301 & ~new_n8092_;
  assign new_n15365_ = ~new_n15363_ & ~new_n15364_;
  assign li0301 = ~lo0055 & ~new_n15365_;
  assign new_n15367_ = lo0937 & new_n4223_;
  assign new_n15368_ = pi059 & ~new_n4223_;
  assign new_n15369_ = ~new_n15367_ & ~new_n15368_;
  assign new_n15370_ = lo0273 & new_n4228_;
  assign new_n15371_ = lo0237 & new_n4219_;
  assign new_n15372_ = ~new_n15370_ & ~new_n15371_;
  assign new_n15373_ = ~new_n4218_ & ~new_n15369_;
  assign li0302 = ~new_n15372_ | new_n15373_;
  assign new_n15375_ = ~lo0478 & lo1043;
  assign new_n15376_ = lo0303 & ~lo1043;
  assign li0303 = new_n15375_ | new_n15376_;
  assign new_n15378_ = ~lo0478 & lo1042;
  assign new_n15379_ = lo0304 & ~lo1042;
  assign li0304 = new_n15378_ | new_n15379_;
  assign new_n15381_ = ~lo0478 & lo1078;
  assign new_n15382_ = lo0305 & ~lo1078;
  assign li0305 = new_n15381_ | new_n15382_;
  assign new_n15384_ = ~lo0478 & lo1053;
  assign new_n15385_ = lo0306 & ~lo1053;
  assign li0306 = new_n15384_ | new_n15385_;
  assign new_n15387_ = ~lo0478 & lo1047;
  assign new_n15388_ = lo0307 & ~lo1047;
  assign li0307 = new_n15387_ | new_n15388_;
  assign new_n15390_ = ~lo0478 & lo1031;
  assign new_n15391_ = lo0308 & ~lo1031;
  assign li0308 = new_n15390_ | new_n15391_;
  assign new_n15393_ = ~lo0478 & lo1066;
  assign new_n15394_ = lo0309 & ~lo1066;
  assign li0309 = new_n15393_ | new_n15394_;
  assign new_n15396_ = lo0934 & new_n4223_;
  assign new_n15397_ = pi058 & ~new_n4223_;
  assign new_n15398_ = ~new_n15396_ & ~new_n15397_;
  assign new_n15399_ = lo0271 & new_n4228_;
  assign new_n15400_ = lo0233 & new_n4219_;
  assign new_n15401_ = ~new_n15399_ & ~new_n15400_;
  assign new_n15402_ = ~new_n4218_ & ~new_n15398_;
  assign li0310 = ~new_n15401_ | new_n15402_;
  assign new_n15404_ = lo0311 & ~new_n8092_;
  assign new_n15405_ = ~lo0311 & ~new_n15360_;
  assign new_n15406_ = lo0311 & new_n15360_;
  assign new_n15407_ = ~new_n15405_ & ~new_n15406_;
  assign new_n15408_ = new_n8092_ & new_n15407_;
  assign new_n15409_ = ~new_n15404_ & ~new_n15408_;
  assign li0311 = ~lo0055 & ~new_n15409_;
  assign new_n15411_ = ~lo0312 & ~new_n8092_;
  assign new_n15412_ = lo0312 & new_n8092_;
  assign new_n15413_ = ~new_n15411_ & ~new_n15412_;
  assign li0312 = ~lo0055 & new_n15413_;
  assign new_n15415_ = lo0314 & li0583;
  assign new_n15416_ = ~new_n4001_ & ~new_n15415_;
  assign new_n15417_ = ~li0583 & ~new_n3985_;
  assign new_n15418_ = new_n3985_ & new_n15416_;
  assign new_n15419_ = new_n4001_ & new_n15417_;
  assign li0477 = ~new_n15418_ & ~new_n15419_;
  assign new_n15421_ = ~lo0954 & ~li0477;
  assign new_n15422_ = lo0313 & lo0954;
  assign li0313 = new_n15421_ | new_n15422_;
  assign new_n15424_ = new_n13252_ & new_n13255_;
  assign new_n15425_ = ~lo0051 & new_n15424_;
  assign new_n15426_ = new_n13236_ & ~new_n13273_;
  assign new_n15427_ = new_n13531_ & new_n15426_;
  assign li0314 = new_n15425_ & new_n15427_;
  assign new_n15429_ = lo0340 & li0480;
  assign new_n15430_ = lo1074 & ~new_n15429_;
  assign new_n15431_ = lo0315 & ~lo1074;
  assign li0315 = new_n15430_ | new_n15431_;
  assign new_n15433_ = lo1041 & ~new_n15429_;
  assign new_n15434_ = lo0316 & ~lo1041;
  assign li0316 = new_n15433_ | new_n15434_;
  assign new_n15436_ = lo0330 & li0480;
  assign new_n15437_ = lo1072 & ~new_n15436_;
  assign new_n15438_ = lo0317 & ~lo1072;
  assign li0317 = new_n15437_ | new_n15438_;
  assign new_n15440_ = lo0341 & li0480;
  assign new_n15441_ = lo1068 & ~new_n15440_;
  assign new_n15442_ = lo0318 & ~lo1068;
  assign li0318 = new_n15441_ | new_n15442_;
  assign new_n15444_ = lo1066 & ~new_n15440_;
  assign new_n15445_ = lo0319 & ~lo1066;
  assign li0319 = new_n15444_ | new_n15445_;
  assign new_n15447_ = lo1042 & ~new_n15429_;
  assign new_n15448_ = lo0320 & ~lo1042;
  assign li0320 = new_n15447_ | new_n15448_;
  assign new_n15450_ = lo1052 & ~new_n15429_;
  assign new_n15451_ = lo0321 & ~lo1052;
  assign li0321 = new_n15450_ | new_n15451_;
  assign new_n15453_ = lo1045 & ~new_n15429_;
  assign new_n15454_ = lo0322 & ~lo1045;
  assign li0322 = new_n15453_ | new_n15454_;
  assign new_n15456_ = lo1059 & ~new_n15429_;
  assign new_n15457_ = lo0323 & ~lo1059;
  assign li0323 = new_n15456_ | new_n15457_;
  assign new_n15459_ = lo1080 & ~new_n15440_;
  assign new_n15460_ = lo0324 & ~lo1080;
  assign li0324 = new_n15459_ | new_n15460_;
  assign new_n15462_ = lo1057 & ~new_n15440_;
  assign new_n15463_ = lo0325 & ~lo1057;
  assign li0325 = new_n15462_ | new_n15463_;
  assign new_n15465_ = lo1051 & ~new_n15440_;
  assign new_n15466_ = lo0326 & ~lo1051;
  assign li0326 = new_n15465_ | new_n15466_;
  assign new_n15468_ = lo1034 & ~new_n15429_;
  assign new_n15469_ = lo0327 & ~lo1034;
  assign li0327 = new_n15468_ | new_n15469_;
  assign new_n15471_ = lo1052 & ~new_n15440_;
  assign new_n15472_ = lo0328 & ~lo1052;
  assign li0328 = new_n15471_ | new_n15472_;
  assign new_n15474_ = lo1037 & ~new_n15440_;
  assign new_n15475_ = lo0329 & ~lo1037;
  assign li0329 = new_n15474_ | new_n15475_;
  assign new_n15477_ = lo0330 & ~li0480;
  assign new_n15478_ = pi003 & ~new_n4666_;
  assign new_n15479_ = ~new_n15429_ & ~new_n15477_;
  assign li0330 = new_n15478_ & ~new_n15479_;
  assign new_n15481_ = lo0331 & ~li0480;
  assign new_n15482_ = ~new_n15440_ & ~new_n15481_;
  assign li0331 = new_n15478_ & ~new_n15482_;
  assign new_n15484_ = ~new_n3628_ & ~new_n3630_;
  assign li0332 = new_n3614_ | ~new_n15484_;
  assign new_n15486_ = lo1034 & ~new_n15440_;
  assign new_n15487_ = lo0333 & ~lo1034;
  assign li0333 = new_n15486_ | new_n15487_;
  assign new_n15489_ = lo1059 & ~new_n15440_;
  assign new_n15490_ = lo0334 & ~lo1059;
  assign li0334 = new_n15489_ | new_n15490_;
  assign new_n15492_ = lo1063 & ~new_n15440_;
  assign new_n15493_ = lo0335 & ~lo1063;
  assign li0335 = new_n15492_ | new_n15493_;
  assign new_n15495_ = lo1064 & ~new_n15436_;
  assign new_n15496_ = lo0336 & ~lo1064;
  assign li0336 = new_n15495_ | new_n15496_;
  assign new_n15498_ = lo1038 & ~new_n15436_;
  assign new_n15499_ = lo0337 & ~lo1038;
  assign li0337 = new_n15498_ | new_n15499_;
  assign new_n15501_ = lo1066 & ~new_n15436_;
  assign new_n15502_ = lo0338 & ~lo1066;
  assign li0338 = new_n15501_ | new_n15502_;
  assign new_n15504_ = lo1080 & ~new_n15436_;
  assign new_n15505_ = lo0339 & ~lo1080;
  assign li0339 = new_n15504_ | new_n15505_;
  assign new_n15507_ = lo0340 & ~li0480;
  assign new_n15508_ = lo0331 & li0480;
  assign new_n15509_ = new_n15478_ & ~new_n15507_;
  assign li0340 = new_n15508_ | ~new_n15509_;
  assign new_n15511_ = lo0341 & ~li0480;
  assign new_n15512_ = ~new_n15436_ & ~new_n15511_;
  assign li0341 = new_n15478_ & ~new_n15512_;
  assign new_n15514_ = lo1043 & ~new_n15429_;
  assign new_n15515_ = lo0342 & ~lo1043;
  assign li0342 = new_n15514_ | new_n15515_;
  assign new_n15517_ = lo1056 & ~new_n15429_;
  assign new_n15518_ = lo0343 & ~lo1056;
  assign li0343 = new_n15517_ | new_n15518_;
  assign new_n15520_ = lo1063 & ~new_n15429_;
  assign new_n15521_ = lo0344 & ~lo1063;
  assign li0344 = new_n15520_ | new_n15521_;
  assign new_n15523_ = lo1033 & ~new_n15429_;
  assign new_n15524_ = lo0345 & ~lo1033;
  assign li0345 = new_n15523_ | new_n15524_;
  assign new_n15526_ = lo1061 & ~new_n15429_;
  assign new_n15527_ = lo0346 & ~lo1061;
  assign li0346 = new_n15526_ | new_n15527_;
  assign new_n15529_ = lo1049 & ~new_n15429_;
  assign new_n15530_ = lo0347 & ~lo1049;
  assign li0347 = new_n15529_ | new_n15530_;
  assign new_n15532_ = lo1081 & ~new_n15429_;
  assign new_n15533_ = lo0348 & ~lo1081;
  assign li0348 = new_n15532_ | new_n15533_;
  assign new_n15535_ = lo1037 & ~new_n15429_;
  assign new_n15536_ = lo0349 & ~lo1037;
  assign li0349 = new_n15535_ | new_n15536_;
  assign new_n15538_ = lo1029 & ~new_n15429_;
  assign new_n15539_ = lo0350 & ~lo1029;
  assign li0350 = new_n15538_ | new_n15539_;
  assign new_n15541_ = lo1073 & ~new_n15429_;
  assign new_n15542_ = lo0351 & ~lo1073;
  assign li0351 = new_n15541_ | new_n15542_;
  assign new_n15544_ = lo1072 & ~new_n15429_;
  assign new_n15545_ = lo0352 & ~lo1072;
  assign li0352 = new_n15544_ | new_n15545_;
  assign new_n15547_ = lo1057 & ~new_n15429_;
  assign new_n15548_ = lo0353 & ~lo1057;
  assign li0353 = new_n15547_ | new_n15548_;
  assign new_n15550_ = lo1039 & ~new_n15429_;
  assign new_n15551_ = lo0354 & ~lo1039;
  assign li0354 = new_n15550_ | new_n15551_;
  assign new_n15553_ = lo1078 & ~new_n15429_;
  assign new_n15554_ = lo0355 & ~lo1078;
  assign li0355 = new_n15553_ | new_n15554_;
  assign new_n15556_ = lo1075 & ~new_n15429_;
  assign new_n15557_ = lo0356 & ~lo1075;
  assign li0356 = new_n15556_ | new_n15557_;
  assign new_n15559_ = lo1070 & ~new_n15429_;
  assign new_n15560_ = lo0357 & ~lo1070;
  assign li0357 = new_n15559_ | new_n15560_;
  assign new_n15562_ = lo1065 & ~new_n15429_;
  assign new_n15563_ = lo0358 & ~lo1065;
  assign li0358 = new_n15562_ | new_n15563_;
  assign new_n15565_ = lo1062 & ~new_n15429_;
  assign new_n15566_ = lo0359 & ~lo1062;
  assign li0359 = new_n15565_ | new_n15566_;
  assign new_n15568_ = lo1036 & ~new_n15429_;
  assign new_n15569_ = lo0360 & ~lo1036;
  assign li0360 = new_n15568_ | new_n15569_;
  assign new_n15571_ = lo1053 & ~new_n15429_;
  assign new_n15572_ = lo0361 & ~lo1053;
  assign li0361 = new_n15571_ | new_n15572_;
  assign new_n15574_ = lo1064 & ~new_n15429_;
  assign new_n15575_ = lo0362 & ~lo1064;
  assign li0362 = new_n15574_ | new_n15575_;
  assign new_n15577_ = lo1043 & ~new_n15436_;
  assign new_n15578_ = lo0363 & ~lo1043;
  assign li0363 = new_n15577_ | new_n15578_;
  assign new_n15580_ = lo1056 & ~new_n15436_;
  assign new_n15581_ = lo0364 & ~lo1056;
  assign li0364 = new_n15580_ | new_n15581_;
  assign new_n15583_ = lo1059 & ~new_n15436_;
  assign new_n15584_ = lo0365 & ~lo1059;
  assign li0365 = new_n15583_ | new_n15584_;
  assign new_n15586_ = lo1063 & ~new_n15436_;
  assign new_n15587_ = lo0366 & ~lo1063;
  assign li0366 = new_n15586_ | new_n15587_;
  assign new_n15589_ = lo1033 & ~new_n15436_;
  assign new_n15590_ = lo0367 & ~lo1033;
  assign li0367 = new_n15589_ | new_n15590_;
  assign new_n15592_ = lo1061 & ~new_n15436_;
  assign new_n15593_ = lo0368 & ~lo1061;
  assign li0368 = new_n15592_ | new_n15593_;
  assign new_n15595_ = lo1074 & ~new_n15436_;
  assign new_n15596_ = lo0369 & ~lo1074;
  assign li0369 = new_n15595_ | new_n15596_;
  assign new_n15598_ = lo1049 & ~new_n15436_;
  assign new_n15599_ = lo0370 & ~lo1049;
  assign li0370 = new_n15598_ | new_n15599_;
  assign new_n15601_ = lo1045 & ~new_n15436_;
  assign new_n15602_ = lo0371 & ~lo1045;
  assign li0371 = new_n15601_ | new_n15602_;
  assign new_n15604_ = lo1042 & ~new_n15436_;
  assign new_n15605_ = lo0372 & ~lo1042;
  assign li0372 = new_n15604_ | new_n15605_;
  assign new_n15607_ = lo1081 & ~new_n15436_;
  assign new_n15608_ = lo0373 & ~lo1081;
  assign li0373 = new_n15607_ | new_n15608_;
  assign new_n15610_ = lo1029 & ~new_n15436_;
  assign new_n15611_ = lo0374 & ~lo1029;
  assign li0374 = new_n15610_ | new_n15611_;
  assign new_n15613_ = lo1041 & ~new_n15436_;
  assign new_n15614_ = lo0375 & ~lo1041;
  assign li0375 = new_n15613_ | new_n15614_;
  assign new_n15616_ = lo1073 & ~new_n15436_;
  assign new_n15617_ = lo0376 & ~lo1073;
  assign li0376 = new_n15616_ | new_n15617_;
  assign new_n15619_ = lo1068 & ~new_n15436_;
  assign new_n15620_ = lo0377 & ~lo1068;
  assign li0377 = new_n15619_ | new_n15620_;
  assign new_n15622_ = lo1057 & ~new_n15436_;
  assign new_n15623_ = lo0378 & ~lo1057;
  assign li0378 = new_n15622_ | new_n15623_;
  assign new_n15625_ = lo1039 & ~new_n15436_;
  assign new_n15626_ = lo0379 & ~lo1039;
  assign li0379 = new_n15625_ | new_n15626_;
  assign new_n15628_ = lo1078 & ~new_n15436_;
  assign new_n15629_ = lo0380 & ~lo1078;
  assign li0380 = new_n15628_ | new_n15629_;
  assign new_n15631_ = lo1075 & ~new_n15436_;
  assign new_n15632_ = lo0381 & ~lo1075;
  assign li0381 = new_n15631_ | new_n15632_;
  assign new_n15634_ = lo1070 & ~new_n15436_;
  assign new_n15635_ = lo0382 & ~lo1070;
  assign li0382 = new_n15634_ | new_n15635_;
  assign new_n15637_ = lo1065 & ~new_n15436_;
  assign new_n15638_ = lo0383 & ~lo1065;
  assign li0383 = new_n15637_ | new_n15638_;
  assign new_n15640_ = lo1062 & ~new_n15436_;
  assign new_n15641_ = lo0384 & ~lo1062;
  assign li0384 = new_n15640_ | new_n15641_;
  assign new_n15643_ = lo1036 & ~new_n15436_;
  assign new_n15644_ = lo0385 & ~lo1036;
  assign li0385 = new_n15643_ | new_n15644_;
  assign new_n15646_ = lo1053 & ~new_n15436_;
  assign new_n15647_ = lo0386 & ~lo1053;
  assign li0386 = new_n15646_ | new_n15647_;
  assign new_n15649_ = lo1047 & ~new_n15436_;
  assign new_n15650_ = lo0387 & ~lo1047;
  assign li0387 = new_n15649_ | new_n15650_;
  assign new_n15652_ = lo1031 & ~new_n15436_;
  assign new_n15653_ = lo0388 & ~lo1031;
  assign li0388 = new_n15652_ | new_n15653_;
  assign new_n15655_ = lo1030 & ~new_n15436_;
  assign new_n15656_ = lo0389 & ~lo1030;
  assign li0389 = new_n15655_ | new_n15656_;
  assign new_n15658_ = lo1043 & ~new_n15440_;
  assign new_n15659_ = lo0390 & ~lo1043;
  assign li0390 = new_n15658_ | new_n15659_;
  assign new_n15661_ = lo1056 & ~new_n15440_;
  assign new_n15662_ = lo0391 & ~lo1056;
  assign li0391 = new_n15661_ | new_n15662_;
  assign new_n15664_ = lo1033 & ~new_n15440_;
  assign new_n15665_ = lo0392 & ~lo1033;
  assign li0392 = new_n15664_ | new_n15665_;
  assign new_n15667_ = lo1061 & ~new_n15440_;
  assign new_n15668_ = lo0393 & ~lo1061;
  assign li0393 = new_n15667_ | new_n15668_;
  assign new_n15670_ = lo1074 & ~new_n15440_;
  assign new_n15671_ = lo0394 & ~lo1074;
  assign li0394 = new_n15670_ | new_n15671_;
  assign new_n15673_ = lo1049 & ~new_n15440_;
  assign new_n15674_ = lo0395 & ~lo1049;
  assign li0395 = new_n15673_ | new_n15674_;
  assign new_n15676_ = lo1045 & ~new_n15440_;
  assign new_n15677_ = lo0396 & ~lo1045;
  assign li0396 = new_n15676_ | new_n15677_;
  assign new_n15679_ = lo1042 & ~new_n15440_;
  assign new_n15680_ = lo0397 & ~lo1042;
  assign li0397 = new_n15679_ | new_n15680_;
  assign new_n15682_ = lo1081 & ~new_n15440_;
  assign new_n15683_ = lo0398 & ~lo1081;
  assign li0398 = new_n15682_ | new_n15683_;
  assign new_n15685_ = lo1041 & ~new_n15440_;
  assign new_n15686_ = lo0399 & ~lo1041;
  assign li0399 = new_n15685_ | new_n15686_;
  assign new_n15688_ = lo1029 & ~new_n15440_;
  assign new_n15689_ = lo0400 & ~lo1029;
  assign li0400 = new_n15688_ | new_n15689_;
  assign new_n15691_ = lo1073 & ~new_n15440_;
  assign new_n15692_ = lo0401 & ~lo1073;
  assign li0401 = new_n15691_ | new_n15692_;
  assign new_n15694_ = lo1072 & ~new_n15440_;
  assign new_n15695_ = lo0402 & ~lo1072;
  assign li0402 = new_n15694_ | new_n15695_;
  assign new_n15697_ = lo1039 & ~new_n15440_;
  assign new_n15698_ = lo0403 & ~lo1039;
  assign li0403 = new_n15697_ | new_n15698_;
  assign new_n15700_ = lo1078 & ~new_n15440_;
  assign new_n15701_ = lo0404 & ~lo1078;
  assign li0404 = new_n15700_ | new_n15701_;
  assign new_n15703_ = lo1075 & ~new_n15440_;
  assign new_n15704_ = lo0405 & ~lo1075;
  assign li0405 = new_n15703_ | new_n15704_;
  assign new_n15706_ = lo1070 & ~new_n15440_;
  assign new_n15707_ = lo0406 & ~lo1070;
  assign li0406 = new_n15706_ | new_n15707_;
  assign new_n15709_ = lo1065 & ~new_n15440_;
  assign new_n15710_ = lo0407 & ~lo1065;
  assign li0407 = new_n15709_ | new_n15710_;
  assign new_n15712_ = lo1062 & ~new_n15440_;
  assign new_n15713_ = lo0408 & ~lo1062;
  assign li0408 = new_n15712_ | new_n15713_;
  assign new_n15715_ = lo1036 & ~new_n15440_;
  assign new_n15716_ = lo0409 & ~lo1036;
  assign li0409 = new_n15715_ | new_n15716_;
  assign new_n15718_ = lo1053 & ~new_n15440_;
  assign new_n15719_ = lo0410 & ~lo1053;
  assign li0410 = new_n15718_ | new_n15719_;
  assign new_n15721_ = lo1047 & ~new_n15440_;
  assign new_n15722_ = lo0411 & ~lo1047;
  assign li0411 = new_n15721_ | new_n15722_;
  assign new_n15724_ = lo1031 & ~new_n15440_;
  assign new_n15725_ = lo0412 & ~lo1031;
  assign li0412 = new_n15724_ | new_n15725_;
  assign new_n15727_ = lo1030 & ~new_n15440_;
  assign new_n15728_ = lo0413 & ~lo1030;
  assign li0413 = new_n15727_ | new_n15728_;
  assign new_n15730_ = lo1043 & ~new_n15508_;
  assign new_n15731_ = lo0414 & ~lo1043;
  assign li0414 = new_n15730_ | new_n15731_;
  assign new_n15733_ = lo1056 & ~new_n15508_;
  assign new_n15734_ = lo0415 & ~lo1056;
  assign li0415 = new_n15733_ | new_n15734_;
  assign new_n15736_ = lo1063 & ~new_n15508_;
  assign new_n15737_ = lo0416 & ~lo1063;
  assign li0416 = new_n15736_ | new_n15737_;
  assign new_n15739_ = lo1033 & ~new_n15508_;
  assign new_n15740_ = lo0417 & ~lo1033;
  assign li0417 = new_n15739_ | new_n15740_;
  assign new_n15742_ = lo1061 & ~new_n15508_;
  assign new_n15743_ = lo0418 & ~lo1061;
  assign li0418 = new_n15742_ | new_n15743_;
  assign new_n15745_ = lo1074 & ~new_n15508_;
  assign new_n15746_ = lo0419 & ~lo1074;
  assign li0419 = new_n15745_ | new_n15746_;
  assign new_n15748_ = lo1049 & ~new_n15508_;
  assign new_n15749_ = lo0420 & ~lo1049;
  assign li0420 = new_n15748_ | new_n15749_;
  assign new_n15751_ = lo1045 & ~new_n15508_;
  assign new_n15752_ = lo0421 & ~lo1045;
  assign li0421 = new_n15751_ | new_n15752_;
  assign new_n15754_ = lo1042 & ~new_n15508_;
  assign new_n15755_ = lo0422 & ~lo1042;
  assign li0422 = new_n15754_ | new_n15755_;
  assign new_n15757_ = lo1081 & ~new_n15508_;
  assign new_n15758_ = lo0423 & ~lo1081;
  assign li0423 = new_n15757_ | new_n15758_;
  assign new_n15760_ = lo1041 & ~new_n15508_;
  assign new_n15761_ = lo0424 & ~lo1041;
  assign li0424 = new_n15760_ | new_n15761_;
  assign new_n15763_ = lo1029 & ~new_n15508_;
  assign new_n15764_ = lo0425 & ~lo1029;
  assign li0425 = new_n15763_ | new_n15764_;
  assign new_n15766_ = lo1073 & ~new_n15508_;
  assign new_n15767_ = lo0426 & ~lo1073;
  assign li0426 = new_n15766_ | new_n15767_;
  assign new_n15769_ = lo1072 & ~new_n15508_;
  assign new_n15770_ = lo0427 & ~lo1072;
  assign li0427 = new_n15769_ | new_n15770_;
  assign new_n15772_ = lo1039 & ~new_n15508_;
  assign new_n15773_ = lo0428 & ~lo1039;
  assign li0428 = new_n15772_ | new_n15773_;
  assign new_n15775_ = lo1078 & ~new_n15508_;
  assign new_n15776_ = lo0429 & ~lo1078;
  assign li0429 = new_n15775_ | new_n15776_;
  assign new_n15778_ = lo1070 & ~new_n15508_;
  assign new_n15779_ = lo0430 & ~lo1070;
  assign li0430 = new_n15778_ | new_n15779_;
  assign new_n15781_ = lo1065 & ~new_n15508_;
  assign new_n15782_ = lo0431 & ~lo1065;
  assign li0431 = new_n15781_ | new_n15782_;
  assign new_n15784_ = lo1062 & ~new_n15508_;
  assign new_n15785_ = lo0432 & ~lo1062;
  assign li0432 = new_n15784_ | new_n15785_;
  assign new_n15787_ = lo1036 & ~new_n15508_;
  assign new_n15788_ = lo0433 & ~lo1036;
  assign li0433 = new_n15787_ | new_n15788_;
  assign new_n15790_ = lo1053 & ~new_n15508_;
  assign new_n15791_ = lo0434 & ~lo1053;
  assign li0434 = new_n15790_ | new_n15791_;
  assign new_n15793_ = lo1047 & ~new_n15508_;
  assign new_n15794_ = lo0435 & ~lo1047;
  assign li0435 = new_n15793_ | new_n15794_;
  assign new_n15796_ = lo1031 & ~new_n15508_;
  assign new_n15797_ = lo0436 & ~lo1031;
  assign li0436 = new_n15796_ | new_n15797_;
  assign new_n15799_ = lo1064 & ~new_n15508_;
  assign new_n15800_ = lo0437 & ~lo1064;
  assign li0437 = new_n15799_ | new_n15800_;
  assign new_n15802_ = lo1030 & ~new_n15508_;
  assign new_n15803_ = lo0438 & ~lo1030;
  assign li0438 = new_n15802_ | new_n15803_;
  assign new_n15805_ = lo1051 & ~new_n15436_;
  assign new_n15806_ = lo0439 & ~lo1051;
  assign li0439 = new_n15805_ | new_n15806_;
  assign new_n15808_ = lo1037 & ~new_n15436_;
  assign new_n15809_ = lo0440 & ~lo1037;
  assign li0440 = new_n15808_ | new_n15809_;
  assign new_n15811_ = lo1038 & ~new_n15429_;
  assign new_n15812_ = lo0441 & ~lo1038;
  assign li0441 = new_n15811_ | new_n15812_;
  assign new_n15814_ = lo1052 & ~new_n15436_;
  assign new_n15815_ = lo0442 & ~lo1052;
  assign li0442 = new_n15814_ | new_n15815_;
  assign new_n15817_ = lo1038 & ~new_n15508_;
  assign new_n15818_ = lo0443 & ~lo1038;
  assign li0443 = new_n15817_ | new_n15818_;
  assign new_n15820_ = lo1066 & ~new_n15508_;
  assign new_n15821_ = lo0444 & ~lo1066;
  assign li0444 = new_n15820_ | new_n15821_;
  assign new_n15823_ = lo1075 & ~new_n15508_;
  assign new_n15824_ = lo0445 & ~lo1075;
  assign li0445 = new_n15823_ | new_n15824_;
  assign new_n15826_ = lo1080 & ~new_n15508_;
  assign new_n15827_ = lo0446 & ~lo1080;
  assign li0446 = new_n15826_ | new_n15827_;
  assign new_n15829_ = lo1034 & ~new_n15436_;
  assign new_n15830_ = lo0447 & ~lo1034;
  assign li0447 = new_n15829_ | new_n15830_;
  assign new_n15832_ = lo1068 & ~new_n15508_;
  assign new_n15833_ = lo0448 & ~lo1068;
  assign li0448 = new_n15832_ | new_n15833_;
  assign new_n15835_ = lo1051 & ~new_n15508_;
  assign new_n15836_ = lo0449 & ~lo1051;
  assign li0449 = new_n15835_ | new_n15836_;
  assign new_n15838_ = lo1030 & ~new_n15429_;
  assign new_n15839_ = lo0450 & ~lo1030;
  assign li0450 = new_n15838_ | new_n15839_;
  assign new_n15841_ = lo1057 & ~new_n15508_;
  assign new_n15842_ = lo0451 & ~lo1057;
  assign li0451 = new_n15841_ | new_n15842_;
  assign new_n15844_ = lo1047 & ~new_n15429_;
  assign new_n15845_ = lo0452 & ~lo1047;
  assign li0452 = new_n15844_ | new_n15845_;
  assign new_n15847_ = lo1034 & ~new_n15508_;
  assign new_n15848_ = lo0453 & ~lo1034;
  assign li0453 = new_n15847_ | new_n15848_;
  assign new_n15850_ = lo1037 & ~new_n15508_;
  assign new_n15851_ = lo0454 & ~lo1037;
  assign li0454 = new_n15850_ | new_n15851_;
  assign new_n15853_ = lo1031 & ~new_n15429_;
  assign new_n15854_ = lo0455 & ~lo1031;
  assign li0455 = new_n15853_ | new_n15854_;
  assign new_n15856_ = lo1038 & ~new_n15440_;
  assign new_n15857_ = lo0456 & ~lo1038;
  assign li0456 = new_n15856_ | new_n15857_;
  assign new_n15859_ = lo0605 & lo0821;
  assign new_n15860_ = lo0600 & lo0601;
  assign new_n15861_ = new_n15859_ & new_n15860_;
  assign new_n15862_ = ~lo0815 & new_n15861_;
  assign new_n15863_ = lo0804 & ~lo0810;
  assign new_n15864_ = lo0804 & lo0810;
  assign new_n15865_ = lo0601 & lo0605;
  assign new_n15866_ = lo0600 & new_n15865_;
  assign new_n15867_ = lo0594 & new_n15866_;
  assign new_n15868_ = lo0821 & new_n15864_;
  assign new_n15869_ = ~lo0815 & new_n15868_;
  assign new_n15870_ = new_n15867_ & new_n15869_;
  assign new_n15871_ = ~lo0804 & ~lo0810;
  assign new_n15872_ = lo0594 & lo0597;
  assign new_n15873_ = new_n15861_ & new_n15871_;
  assign new_n15874_ = lo0815 & new_n15873_;
  assign new_n15875_ = new_n15872_ & new_n15874_;
  assign new_n15876_ = ~lo0804 & lo0810;
  assign new_n15877_ = new_n15859_ & new_n15876_;
  assign new_n15878_ = ~lo0815 & new_n15877_;
  assign new_n15879_ = lo0601 & new_n15878_;
  assign new_n15880_ = lo0821 & new_n15860_;
  assign new_n15881_ = lo0605 & new_n15880_;
  assign new_n15882_ = lo0599 & new_n15881_;
  assign new_n15883_ = lo0594 & new_n15882_;
  assign new_n15884_ = lo0597 & new_n15883_;
  assign new_n15885_ = lo0595 & lo0596;
  assign new_n15886_ = new_n15864_ & new_n15884_;
  assign new_n15887_ = lo0815 & new_n15886_;
  assign new_n15888_ = new_n15885_ & new_n15887_;
  assign new_n15889_ = ~new_n15870_ & ~new_n15875_;
  assign new_n15890_ = ~new_n15879_ & new_n15889_;
  assign new_n15891_ = ~new_n15888_ & new_n15890_;
  assign new_n15892_ = new_n15862_ & new_n15863_;
  assign new_n15893_ = new_n15891_ & ~new_n15892_;
  assign new_n15894_ = lo0601 & lo0815;
  assign new_n15895_ = lo0594 & lo0600;
  assign new_n15896_ = new_n15894_ & new_n15895_;
  assign new_n15897_ = lo0595 & lo0597;
  assign new_n15898_ = new_n15876_ & new_n15896_;
  assign new_n15899_ = new_n15897_ & new_n15898_;
  assign new_n15900_ = new_n15859_ & new_n15899_;
  assign new_n15901_ = new_n15880_ & new_n15897_;
  assign new_n15902_ = lo0594 & lo0605;
  assign new_n15903_ = lo0596 & new_n15902_;
  assign new_n15904_ = new_n15901_ & new_n15903_;
  assign new_n15905_ = new_n15863_ & new_n15904_;
  assign new_n15906_ = lo0815 & new_n15905_;
  assign new_n15907_ = new_n15859_ & new_n15871_;
  assign new_n15908_ = ~lo0815 & new_n15907_;
  assign new_n15909_ = new_n15893_ & ~new_n15900_;
  assign new_n15910_ = ~new_n15906_ & new_n15909_;
  assign li0457 = new_n15908_ | ~new_n15910_;
  assign new_n15912_ = lo1066 & ~new_n15429_;
  assign new_n15913_ = lo0458 & ~lo1066;
  assign li0458 = new_n15912_ | new_n15913_;
  assign new_n15915_ = lo1052 & ~new_n15508_;
  assign new_n15916_ = lo0459 & ~lo1052;
  assign li0459 = new_n15915_ | new_n15916_;
  assign new_n15918_ = lo1080 & ~new_n15429_;
  assign new_n15919_ = lo0460 & ~lo1080;
  assign li0460 = new_n15918_ | new_n15919_;
  assign new_n15921_ = lo1051 & ~new_n15429_;
  assign new_n15922_ = lo0461 & ~lo1051;
  assign li0461 = new_n15921_ | new_n15922_;
  assign new_n15924_ = lo1068 & ~new_n15429_;
  assign new_n15925_ = lo0462 & ~lo1068;
  assign li0462 = new_n15924_ | new_n15925_;
  assign new_n15927_ = lo1064 & ~new_n15440_;
  assign new_n15928_ = lo0463 & ~lo1064;
  assign li0463 = new_n15927_ | new_n15928_;
  assign new_n15930_ = lo1059 & ~new_n15508_;
  assign new_n15931_ = lo0464 & ~lo1059;
  assign li0464 = new_n15930_ | new_n15931_;
  assign new_n15933_ = lo0926 & new_n4223_;
  assign new_n15934_ = pi068 & ~new_n4223_;
  assign new_n15935_ = ~new_n15933_ & ~new_n15934_;
  assign new_n15936_ = ~new_n4218_ & ~new_n15935_;
  assign new_n15937_ = lo0243 & new_n4228_;
  assign li0465 = new_n15936_ | new_n15937_;
  assign new_n15939_ = lo0943 & new_n4223_;
  assign new_n15940_ = pi062 & ~new_n4223_;
  assign new_n15941_ = ~new_n15939_ & ~new_n15940_;
  assign new_n15942_ = ~new_n4218_ & ~new_n15941_;
  assign new_n15943_ = lo0275 & new_n4228_;
  assign li0466 = new_n15942_ | new_n15943_;
  assign new_n15945_ = ~lo0995 & new_n4524_;
  assign new_n15946_ = lo0040 & li0793;
  assign new_n15947_ = new_n4167_ & new_n4175_;
  assign new_n15948_ = ~lo0040 & new_n3548_;
  assign new_n15949_ = new_n4170_ & new_n15947_;
  assign new_n15950_ = new_n4185_ & new_n15949_;
  assign new_n15951_ = new_n15948_ & new_n15950_;
  assign new_n15952_ = new_n4176_ & new_n14230_;
  assign new_n15953_ = new_n15951_ & new_n15952_;
  assign new_n15954_ = new_n4189_ & new_n15953_;
  assign new_n15955_ = new_n3549_ & new_n15954_;
  assign new_n15956_ = new_n4171_ & new_n15955_;
  assign new_n15957_ = lo0065 & lo0102;
  assign new_n15958_ = ~lo0065 & ~lo0102;
  assign new_n15959_ = ~new_n15957_ & ~new_n15958_;
  assign new_n15960_ = new_n15956_ & new_n15959_;
  assign new_n15961_ = ~lo0048 & new_n4194_;
  assign new_n15962_ = new_n4153_ & new_n4154_;
  assign new_n15963_ = new_n15960_ & new_n15962_;
  assign new_n15964_ = new_n15961_ & new_n15963_;
  assign new_n15965_ = new_n13344_ & new_n15964_;
  assign new_n15966_ = ~lo0040 & new_n15965_;
  assign new_n15967_ = ~li0893 & new_n15966_;
  assign new_n15968_ = new_n13357_ & new_n13363_;
  assign new_n15969_ = new_n15967_ & new_n15968_;
  assign new_n15970_ = ~lo0984 & new_n15946_;
  assign new_n15971_ = new_n15945_ & new_n15970_;
  assign li0467 = new_n15969_ | new_n15971_;
  assign new_n15973_ = lo0024 & new_n3618_;
  assign new_n15974_ = new_n4525_ & new_n7791_;
  assign new_n15975_ = lo0468 & ~new_n15973_;
  assign li0468 = new_n15974_ | new_n15975_;
  assign new_n15977_ = lo0942 & new_n4223_;
  assign new_n15978_ = pi067 & ~new_n4223_;
  assign new_n15979_ = ~new_n15977_ & ~new_n15978_;
  assign new_n15980_ = ~new_n4218_ & ~new_n15979_;
  assign new_n15981_ = lo0263 & new_n4228_;
  assign li0469 = new_n15980_ | new_n15981_;
  assign new_n15983_ = lo0925 & new_n4223_;
  assign new_n15984_ = pi066 & ~new_n4223_;
  assign new_n15985_ = ~new_n15983_ & ~new_n15984_;
  assign new_n15986_ = ~new_n4218_ & ~new_n15985_;
  assign new_n15987_ = lo0267 & new_n4228_;
  assign li0470 = new_n15986_ | new_n15987_;
  assign new_n15989_ = lo0941 & new_n4223_;
  assign new_n15990_ = pi064 & ~new_n4223_;
  assign new_n15991_ = ~new_n15989_ & ~new_n15990_;
  assign new_n15992_ = ~new_n4218_ & ~new_n15991_;
  assign new_n15993_ = lo0253 & new_n4228_;
  assign li0471 = new_n15992_ | new_n15993_;
  assign new_n15995_ = lo0923 & new_n4223_;
  assign new_n15996_ = pi065 & ~new_n4223_;
  assign new_n15997_ = ~new_n15995_ & ~new_n15996_;
  assign new_n15998_ = ~new_n4218_ & ~new_n15997_;
  assign new_n15999_ = lo0254 & new_n4228_;
  assign li0472 = new_n15998_ | new_n15999_;
  assign new_n16001_ = lo0922 & new_n4223_;
  assign new_n16002_ = pi063 & ~new_n4223_;
  assign new_n16003_ = ~new_n16001_ & ~new_n16002_;
  assign new_n16004_ = ~new_n4218_ & ~new_n16003_;
  assign new_n16005_ = lo0268 & new_n4228_;
  assign li0473 = new_n16004_ | new_n16005_;
  assign new_n16007_ = lo0931 & new_n4223_;
  assign new_n16008_ = pi061 & ~new_n4223_;
  assign new_n16009_ = ~new_n16007_ & ~new_n16008_;
  assign new_n16010_ = ~new_n4218_ & ~new_n16009_;
  assign new_n16011_ = lo0272 & new_n4228_;
  assign li0474 = new_n16010_ | new_n16011_;
  assign new_n16013_ = lo0936 & new_n4223_;
  assign new_n16014_ = pi060 & ~new_n4223_;
  assign new_n16015_ = ~new_n16013_ & ~new_n16014_;
  assign new_n16016_ = ~new_n4218_ & ~new_n16015_;
  assign new_n16017_ = lo0283 & new_n4228_;
  assign li0475 = new_n16016_ | new_n16017_;
  assign new_n16019_ = ~lo0060 & ~lo0061;
  assign new_n16020_ = new_n13362_ & new_n16019_;
  assign new_n16021_ = new_n13344_ & new_n16020_;
  assign new_n16022_ = new_n15338_ & new_n16021_;
  assign new_n16023_ = new_n4158_ & new_n5297_;
  assign new_n16024_ = new_n16022_ & new_n16023_;
  assign new_n16025_ = new_n4185_ & new_n13354_;
  assign new_n16026_ = new_n4189_ & new_n16025_;
  assign new_n16027_ = ~lo0048 & new_n16026_;
  assign new_n16028_ = lo0084 & new_n16027_;
  assign new_n16029_ = new_n4174_ & new_n16028_;
  assign new_n16030_ = new_n16024_ & new_n16029_;
  assign new_n16031_ = new_n13355_ & new_n16030_;
  assign new_n16032_ = new_n4194_ & new_n16031_;
  assign new_n16033_ = ~lo0051 & ~lo0081;
  assign new_n16034_ = new_n4177_ & new_n13346_;
  assign new_n16035_ = new_n3557_ & new_n16034_;
  assign new_n16036_ = new_n16033_ & new_n16035_;
  assign new_n16037_ = ~li0893 & new_n16036_;
  assign new_n16038_ = ~lo0071 & new_n16037_;
  assign new_n16039_ = ~lo0046 & new_n16038_;
  assign new_n16040_ = ~lo0068 & new_n16039_;
  assign new_n16041_ = lo0071 & new_n8536_;
  assign new_n16042_ = new_n16032_ & new_n16040_;
  assign li0476 = new_n16041_ | new_n16042_;
  assign li0478 = lo0071 & new_n6074_;
  assign new_n16045_ = lo0248 & ~new_n14275_;
  assign new_n16046_ = ~lo0248 & lo0481;
  assign li0481 = new_n16045_ | new_n16046_;
  assign new_n16048_ = lo0249 & ~new_n14289_;
  assign new_n16049_ = ~lo0249 & lo0482;
  assign li0482 = new_n16048_ | new_n16049_;
  assign new_n16051_ = lo0242 & ~new_n14310_;
  assign new_n16052_ = ~lo0242 & lo0483;
  assign li0483 = new_n16051_ | new_n16052_;
  assign new_n16054_ = lo0249 & ~new_n14310_;
  assign new_n16055_ = ~lo0249 & lo0484;
  assign li0484 = new_n16054_ | new_n16055_;
  assign new_n16057_ = lo0234 & ~new_n14386_;
  assign new_n16058_ = ~lo0234 & lo0485;
  assign li0485 = new_n16057_ | new_n16058_;
  assign new_n16060_ = lo0244 & ~new_n14386_;
  assign new_n16061_ = ~lo0244 & lo0486;
  assign li0486 = new_n16060_ | new_n16061_;
  assign new_n16063_ = lo0246 & ~new_n14275_;
  assign new_n16064_ = ~lo0246 & lo0487;
  assign li0487 = new_n16063_ | new_n16064_;
  assign new_n16066_ = lo0239 & ~new_n14275_;
  assign new_n16067_ = ~lo0239 & lo0488;
  assign li0488 = new_n16066_ | new_n16067_;
  assign new_n16069_ = lo0242 & ~new_n14386_;
  assign new_n16070_ = ~lo0242 & lo0489;
  assign li0489 = new_n16069_ | new_n16070_;
  assign new_n16072_ = lo0241 & ~new_n14310_;
  assign new_n16073_ = ~lo0241 & lo0490;
  assign li0490 = new_n16072_ | new_n16073_;
  assign new_n16075_ = lo0238 & ~new_n14310_;
  assign new_n16076_ = ~lo0238 & lo0491;
  assign li0491 = new_n16075_ | new_n16076_;
  assign new_n16078_ = lo0240 & ~new_n14310_;
  assign new_n16079_ = ~lo0240 & lo0492;
  assign li0492 = new_n16078_ | new_n16079_;
  assign new_n16081_ = lo0244 & ~new_n14310_;
  assign new_n16082_ = ~lo0244 & lo0493;
  assign li0493 = new_n16081_ | new_n16082_;
  assign new_n16084_ = lo0239 & ~new_n14310_;
  assign new_n16085_ = ~lo0239 & lo0494;
  assign li0494 = new_n16084_ | new_n16085_;
  assign new_n16087_ = lo0235 & ~new_n14310_;
  assign new_n16088_ = ~lo0235 & lo0495;
  assign li0495 = new_n16087_ | new_n16088_;
  assign new_n16090_ = lo0249 & ~new_n14304_;
  assign new_n16091_ = ~lo0249 & lo0496;
  assign li0496 = new_n16090_ | new_n16091_;
  assign new_n16093_ = lo0239 & ~new_n14304_;
  assign new_n16094_ = ~lo0239 & lo0497;
  assign li0497 = new_n16093_ | new_n16094_;
  assign new_n16096_ = lo0238 & ~new_n14289_;
  assign new_n16097_ = ~lo0238 & lo0498;
  assign li0498 = new_n16096_ | new_n16097_;
  assign new_n16099_ = lo0246 & ~new_n14304_;
  assign new_n16100_ = ~lo0246 & lo0499;
  assign li0499 = new_n16099_ | new_n16100_;
  assign new_n16102_ = lo0241 & ~new_n14304_;
  assign new_n16103_ = ~lo0241 & lo0500;
  assign li0500 = new_n16102_ | new_n16103_;
  assign new_n16105_ = lo0248 & ~new_n14304_;
  assign new_n16106_ = ~lo0248 & lo0501;
  assign li0501 = new_n16105_ | new_n16106_;
  assign new_n16108_ = lo0247 & ~new_n14304_;
  assign new_n16109_ = ~lo0247 & lo0502;
  assign li0502 = new_n16108_ | new_n16109_;
  assign new_n16111_ = lo0245 & ~new_n14304_;
  assign new_n16112_ = ~lo0245 & lo0503;
  assign li0503 = new_n16111_ | new_n16112_;
  assign new_n16114_ = lo0242 & ~new_n14297_;
  assign new_n16115_ = ~lo0242 & lo0504;
  assign li0504 = new_n16114_ | new_n16115_;
  assign new_n16117_ = lo0234 & ~new_n14304_;
  assign new_n16118_ = ~lo0234 & lo0505;
  assign li0505 = new_n16117_ | new_n16118_;
  assign new_n16120_ = lo0241 & ~new_n14297_;
  assign new_n16121_ = ~lo0241 & lo0506;
  assign li0506 = new_n16120_ | new_n16121_;
  assign new_n16123_ = lo0238 & ~new_n14297_;
  assign new_n16124_ = ~lo0238 & lo0507;
  assign li0507 = new_n16123_ | new_n16124_;
  assign new_n16126_ = lo0247 & ~new_n14297_;
  assign new_n16127_ = ~lo0247 & lo0508;
  assign li0508 = new_n16126_ | new_n16127_;
  assign new_n16129_ = lo0245 & ~new_n14297_;
  assign new_n16130_ = ~lo0245 & lo0509;
  assign li0509 = new_n16129_ | new_n16130_;
  assign new_n16132_ = lo0242 & ~new_n14275_;
  assign new_n16133_ = ~lo0242 & lo0510;
  assign li0510 = new_n16132_ | new_n16133_;
  assign new_n16135_ = lo0234 & ~new_n14275_;
  assign new_n16136_ = ~lo0234 & lo0511;
  assign li0511 = new_n16135_ | new_n16136_;
  assign new_n16138_ = lo0235 & ~new_n14275_;
  assign new_n16139_ = ~lo0235 & lo0512;
  assign li0512 = new_n16138_ | new_n16139_;
  assign new_n16141_ = lo0244 & ~new_n14275_;
  assign new_n16142_ = ~lo0244 & lo0513;
  assign li0513 = new_n16141_ | new_n16142_;
  assign new_n16144_ = lo0245 & ~new_n14275_;
  assign new_n16145_ = ~lo0245 & lo0514;
  assign li0514 = new_n16144_ | new_n16145_;
  assign new_n16147_ = lo0240 & ~new_n14275_;
  assign new_n16148_ = ~lo0240 & lo0515;
  assign li0515 = new_n16147_ | new_n16148_;
  assign new_n16150_ = lo0247 & ~new_n14275_;
  assign new_n16151_ = ~lo0247 & lo0516;
  assign li0516 = new_n16150_ | new_n16151_;
  assign new_n16153_ = lo0238 & ~new_n14275_;
  assign new_n16154_ = ~lo0238 & lo0517;
  assign li0517 = new_n16153_ | new_n16154_;
  assign new_n16156_ = lo0234 & ~new_n14283_;
  assign new_n16157_ = ~lo0234 & lo0518;
  assign li0518 = new_n16156_ | new_n16157_;
  assign new_n16159_ = lo0239 & ~new_n14283_;
  assign new_n16160_ = ~lo0239 & lo0519;
  assign li0519 = new_n16159_ | new_n16160_;
  assign new_n16162_ = lo0246 & ~new_n14283_;
  assign new_n16163_ = ~lo0246 & lo0520;
  assign li0520 = new_n16162_ | new_n16163_;
  assign new_n16165_ = lo0248 & ~new_n14283_;
  assign new_n16166_ = ~lo0248 & lo0521;
  assign li0521 = new_n16165_ | new_n16166_;
  assign new_n16168_ = lo0238 & ~new_n14283_;
  assign new_n16169_ = ~lo0238 & lo0522;
  assign li0522 = new_n16168_ | new_n16169_;
  assign new_n16171_ = lo0234 & ~new_n14397_;
  assign new_n16172_ = ~lo0234 & lo0523;
  assign li0523 = new_n16171_ | new_n16172_;
  assign new_n16174_ = lo0239 & ~new_n14397_;
  assign new_n16175_ = ~lo0239 & lo0524;
  assign li0524 = new_n16174_ | new_n16175_;
  assign new_n16177_ = lo0245 & ~new_n14397_;
  assign new_n16178_ = ~lo0245 & lo0525;
  assign li0525 = new_n16177_ | new_n16178_;
  assign new_n16180_ = lo0246 & ~new_n14397_;
  assign new_n16181_ = ~lo0246 & lo0526;
  assign li0526 = new_n16180_ | new_n16181_;
  assign new_n16183_ = lo0247 & ~new_n14397_;
  assign new_n16184_ = ~lo0247 & lo0527;
  assign li0527 = new_n16183_ | new_n16184_;
  assign new_n16186_ = lo0249 & ~new_n14397_;
  assign new_n16187_ = ~lo0249 & lo0528;
  assign li0528 = new_n16186_ | new_n16187_;
  assign new_n16189_ = lo0238 & ~new_n14397_;
  assign new_n16190_ = ~lo0238 & lo0529;
  assign li0529 = new_n16189_ | new_n16190_;
  assign new_n16192_ = lo0240 & ~new_n14397_;
  assign new_n16193_ = ~lo0240 & lo0530;
  assign li0530 = new_n16192_ | new_n16193_;
  assign new_n16195_ = lo0235 & ~new_n14289_;
  assign new_n16196_ = ~lo0235 & lo0531;
  assign li0531 = new_n16195_ | new_n16196_;
  assign new_n16198_ = lo0247 & ~new_n14289_;
  assign new_n16199_ = ~lo0247 & lo0532;
  assign li0532 = new_n16198_ | new_n16199_;
  assign new_n16201_ = lo0235 & ~new_n14297_;
  assign new_n16202_ = ~lo0235 & lo0533;
  assign li0533 = new_n16201_ | new_n16202_;
  assign new_n16204_ = lo0239 & ~new_n14297_;
  assign new_n16205_ = ~lo0239 & lo0534;
  assign li0534 = new_n16204_ | new_n16205_;
  assign new_n16207_ = lo0240 & ~new_n14297_;
  assign new_n16208_ = ~lo0240 & lo0535;
  assign li0535 = new_n16207_ | new_n16208_;
  assign new_n16210_ = lo0246 & ~new_n14297_;
  assign new_n16211_ = ~lo0246 & lo0536;
  assign li0536 = new_n16210_ | new_n16211_;
  assign new_n16213_ = lo0248 & ~new_n14297_;
  assign new_n16214_ = ~lo0248 & lo0537;
  assign li0537 = new_n16213_ | new_n16214_;
  assign new_n16216_ = lo0249 & ~new_n14297_;
  assign new_n16217_ = ~lo0249 & lo0538;
  assign li0538 = new_n16216_ | new_n16217_;
  assign new_n16219_ = lo0242 & ~new_n14304_;
  assign new_n16220_ = ~lo0242 & lo0539;
  assign li0539 = new_n16219_ | new_n16220_;
  assign new_n16222_ = lo0235 & ~new_n14304_;
  assign new_n16223_ = ~lo0235 & lo0540;
  assign li0540 = new_n16222_ | new_n16223_;
  assign new_n16225_ = lo0244 & ~new_n14304_;
  assign new_n16226_ = ~lo0244 & lo0541;
  assign li0541 = new_n16225_ | new_n16226_;
  assign new_n16228_ = lo0240 & ~new_n14304_;
  assign new_n16229_ = ~lo0240 & lo0542;
  assign li0542 = new_n16228_ | new_n16229_;
  assign new_n16231_ = lo0238 & ~new_n14304_;
  assign new_n16232_ = ~lo0238 & lo0543;
  assign li0543 = new_n16231_ | new_n16232_;
  assign new_n16234_ = lo0234 & ~new_n14310_;
  assign new_n16235_ = ~lo0234 & lo0544;
  assign li0544 = new_n16234_ | new_n16235_;
  assign new_n16237_ = lo0245 & ~new_n14310_;
  assign new_n16238_ = ~lo0245 & lo0545;
  assign li0545 = new_n16237_ | new_n16238_;
  assign new_n16240_ = lo0246 & ~new_n14310_;
  assign new_n16241_ = ~lo0246 & lo0546;
  assign li0546 = new_n16240_ | new_n16241_;
  assign new_n16243_ = lo0247 & ~new_n14310_;
  assign new_n16244_ = ~lo0247 & lo0547;
  assign li0547 = new_n16243_ | new_n16244_;
  assign new_n16246_ = lo0248 & ~new_n14310_;
  assign new_n16247_ = ~lo0248 & lo0548;
  assign li0548 = new_n16246_ | new_n16247_;
  assign new_n16249_ = lo0235 & ~new_n14386_;
  assign new_n16250_ = ~lo0235 & lo0549;
  assign li0549 = new_n16249_ | new_n16250_;
  assign new_n16252_ = lo0239 & ~new_n14386_;
  assign new_n16253_ = ~lo0239 & lo0550;
  assign li0550 = new_n16252_ | new_n16253_;
  assign new_n16255_ = lo0240 & ~new_n14386_;
  assign new_n16256_ = ~lo0240 & lo0551;
  assign li0551 = new_n16255_ | new_n16256_;
  assign new_n16258_ = lo0247 & ~new_n14386_;
  assign new_n16259_ = ~lo0247 & lo0552;
  assign li0552 = new_n16258_ | new_n16259_;
  assign new_n16261_ = lo0241 & ~new_n14386_;
  assign new_n16262_ = ~lo0241 & lo0553;
  assign li0553 = new_n16261_ | new_n16262_;
  assign new_n16264_ = lo0248 & ~new_n14386_;
  assign new_n16265_ = ~lo0248 & lo0554;
  assign li0554 = new_n16264_ | new_n16265_;
  assign new_n16267_ = lo0249 & ~new_n14386_;
  assign new_n16268_ = ~lo0249 & lo0555;
  assign li0555 = new_n16267_ | new_n16268_;
  assign new_n16270_ = lo0242 & ~new_n14289_;
  assign new_n16271_ = ~lo0242 & lo0556;
  assign li0556 = new_n16270_ | new_n16271_;
  assign new_n16273_ = lo0234 & ~new_n14297_;
  assign new_n16274_ = ~lo0234 & lo0557;
  assign li0557 = new_n16273_ | new_n16274_;
  assign new_n16276_ = lo0244 & ~new_n14297_;
  assign new_n16277_ = ~lo0244 & lo0558;
  assign li0558 = new_n16276_ | new_n16277_;
  assign new_n16279_ = lo0241 & ~new_n14275_;
  assign new_n16280_ = ~lo0241 & lo0559;
  assign li0559 = new_n16279_ | new_n16280_;
  assign new_n16282_ = lo0240 & ~new_n14289_;
  assign new_n16283_ = ~lo0240 & lo0560;
  assign li0560 = new_n16282_ | new_n16283_;
  assign new_n16285_ = lo0247 & ~new_n14283_;
  assign new_n16286_ = ~lo0247 & lo0561;
  assign li0561 = new_n16285_ | new_n16286_;
  assign new_n16288_ = lo0241 & ~new_n14289_;
  assign new_n16289_ = ~lo0241 & lo0562;
  assign li0562 = new_n16288_ | new_n16289_;
  assign new_n16291_ = lo0246 & ~new_n14386_;
  assign new_n16292_ = ~lo0246 & lo0563;
  assign li0563 = new_n16291_ | new_n16292_;
  assign new_n16294_ = lo0246 & ~new_n14289_;
  assign new_n16295_ = ~lo0246 & lo0564;
  assign li0564 = new_n16294_ | new_n16295_;
  assign new_n16297_ = lo0248 & ~new_n14289_;
  assign new_n16298_ = ~lo0248 & lo0565;
  assign li0565 = new_n16297_ | new_n16298_;
  assign new_n16300_ = lo0244 & ~new_n14289_;
  assign new_n16301_ = ~lo0244 & lo0566;
  assign li0566 = new_n16300_ | new_n16301_;
  assign li0946 = lo0230 & new_n3673_;
  assign new_n16304_ = lo0567 & ~li0946;
  assign new_n16305_ = pi003 & new_n16304_;
  assign new_n16306_ = lo0665 & new_n13784_;
  assign new_n16307_ = lo0621 & new_n13735_;
  assign new_n16308_ = ~new_n16306_ & ~new_n16307_;
  assign new_n16309_ = li0946 & ~new_n16308_;
  assign new_n16310_ = pi002 & new_n16309_;
  assign li0567 = new_n16305_ | new_n16310_;
  assign new_n16312_ = lo0245 & ~new_n14289_;
  assign new_n16313_ = ~lo0245 & lo0568;
  assign li0568 = new_n16312_ | new_n16313_;
  assign new_n16315_ = lo0239 & ~new_n14289_;
  assign new_n16316_ = ~lo0239 & lo0569;
  assign li0569 = new_n16315_ | new_n16316_;
  assign new_n16318_ = lo0234 & ~new_n14289_;
  assign new_n16319_ = ~lo0234 & lo0570;
  assign li0570 = new_n16318_ | new_n16319_;
  assign new_n16321_ = lo0241 & ~new_n14397_;
  assign new_n16322_ = ~lo0241 & lo0571;
  assign li0571 = new_n16321_ | new_n16322_;
  assign new_n16324_ = lo0244 & ~new_n14397_;
  assign new_n16325_ = ~lo0244 & lo0572;
  assign li0572 = new_n16324_ | new_n16325_;
  assign new_n16327_ = lo0242 & ~new_n14397_;
  assign new_n16328_ = ~lo0242 & lo0573;
  assign li0573 = new_n16327_ | new_n16328_;
  assign new_n16330_ = lo0241 & ~new_n14283_;
  assign new_n16331_ = ~lo0241 & lo0574;
  assign li0574 = new_n16330_ | new_n16331_;
  assign new_n16333_ = lo0235 & ~new_n14397_;
  assign new_n16334_ = ~lo0235 & lo0575;
  assign li0575 = new_n16333_ | new_n16334_;
  assign new_n16336_ = lo0248 & ~new_n14397_;
  assign new_n16337_ = ~lo0248 & lo0576;
  assign li0576 = new_n16336_ | new_n16337_;
  assign new_n16339_ = lo0238 & ~new_n14386_;
  assign new_n16340_ = ~lo0238 & lo0577;
  assign li0577 = new_n16339_ | new_n16340_;
  assign new_n16342_ = lo0249 & ~new_n14283_;
  assign new_n16343_ = ~lo0249 & lo0578;
  assign li0578 = new_n16342_ | new_n16343_;
  assign new_n16345_ = lo0249 & ~new_n14275_;
  assign new_n16346_ = ~lo0249 & lo0579;
  assign li0579 = new_n16345_ | new_n16346_;
  assign new_n16348_ = lo0245 & ~new_n14386_;
  assign new_n16349_ = ~lo0245 & lo0580;
  assign li0580 = new_n16348_ | new_n16349_;
  assign new_n16351_ = lo0235 & ~new_n14283_;
  assign new_n16352_ = ~lo0235 & lo0581;
  assign li0581 = new_n16351_ | new_n16352_;
  assign new_n16354_ = lo0240 & ~new_n14283_;
  assign new_n16355_ = ~lo0240 & lo0582;
  assign li0582 = new_n16354_ | new_n16355_;
  assign new_n16357_ = lo0245 & ~new_n14283_;
  assign new_n16358_ = ~lo0245 & lo0584;
  assign li0584 = new_n16357_ | new_n16358_;
  assign new_n16360_ = lo0244 & ~new_n14283_;
  assign new_n16361_ = ~lo0244 & lo0585;
  assign li0585 = new_n16360_ | new_n16361_;
  assign new_n16363_ = lo0242 & ~new_n14283_;
  assign new_n16364_ = ~lo0242 & lo0586;
  assign li0586 = new_n16363_ | new_n16364_;
  assign new_n16366_ = lo0230 & lo0587;
  assign new_n16367_ = ~lo0587 & new_n13737_;
  assign li0587 = new_n16366_ | new_n16367_;
  assign new_n16369_ = lo0123 & new_n3678_;
  assign new_n16370_ = lo0588 & ~new_n16369_;
  assign new_n16371_ = lo0591 & new_n16369_;
  assign new_n16372_ = ~new_n16370_ & ~new_n16371_;
  assign li0588 = new_n15478_ & ~new_n16372_;
  assign new_n16374_ = lo0201 & new_n14213_;
  assign new_n16375_ = lo0202 & new_n14278_;
  assign new_n16376_ = ~new_n16374_ & ~new_n16375_;
  assign new_n16377_ = lo0220 & new_n14306_;
  assign new_n16378_ = lo0203 & new_n14285_;
  assign new_n16379_ = ~new_n16377_ & ~new_n16378_;
  assign new_n16380_ = new_n16376_ & new_n16379_;
  assign new_n16381_ = new_n4460_ & ~new_n16380_;
  assign new_n16382_ = lo0204 & new_n14213_;
  assign new_n16383_ = lo0205 & new_n14278_;
  assign new_n16384_ = ~new_n16382_ & ~new_n16383_;
  assign new_n16385_ = lo0218 & new_n14285_;
  assign new_n16386_ = new_n16384_ & ~new_n16385_;
  assign new_n16387_ = lo0206 & new_n14306_;
  assign new_n16388_ = new_n16386_ & ~new_n16387_;
  assign new_n16389_ = ~new_n4469_ & ~new_n16388_;
  assign li0589 = new_n16381_ | new_n16389_;
  assign new_n16391_ = lo0588 & new_n16369_;
  assign new_n16392_ = lo0590 & ~new_n16369_;
  assign new_n16393_ = ~new_n16391_ & ~new_n16392_;
  assign li0590 = ~new_n15478_ | ~new_n16393_;
  assign new_n16395_ = lo0591 & ~new_n16369_;
  assign new_n16396_ = lo0592 & new_n16369_;
  assign new_n16397_ = ~new_n16395_ & ~new_n16396_;
  assign li0591 = new_n15478_ & ~new_n16397_;
  assign new_n16399_ = lo0592 & ~new_n16369_;
  assign new_n16400_ = lo0590 & new_n16369_;
  assign new_n16401_ = ~new_n16399_ & ~new_n16400_;
  assign li0592 = new_n15478_ & ~new_n16401_;
  assign new_n16403_ = lo0239 & ~lo0497;
  assign new_n16404_ = ~new_n16094_ & ~new_n16403_;
  assign new_n16405_ = lo0246 & lo0499;
  assign new_n16406_ = ~lo0246 & ~lo0499;
  assign new_n16407_ = ~new_n16405_ & ~new_n16406_;
  assign new_n16408_ = new_n14278_ & ~new_n16407_;
  assign new_n16409_ = lo0248 & ~lo0501;
  assign new_n16410_ = ~new_n16106_ & ~new_n16409_;
  assign new_n16411_ = new_n16408_ & new_n16410_;
  assign new_n16412_ = lo0247 & ~lo0502;
  assign new_n16413_ = ~new_n16109_ & ~new_n16412_;
  assign new_n16414_ = lo0241 & ~lo0500;
  assign new_n16415_ = ~new_n16103_ & ~new_n16414_;
  assign new_n16416_ = new_n16413_ & new_n16415_;
  assign new_n16417_ = lo0235 & ~lo0540;
  assign new_n16418_ = ~new_n16223_ & ~new_n16417_;
  assign new_n16419_ = lo0238 & ~lo0543;
  assign new_n16420_ = ~new_n16232_ & ~new_n16419_;
  assign new_n16421_ = new_n16418_ & new_n16420_;
  assign new_n16422_ = lo0249 & ~lo0496;
  assign new_n16423_ = ~new_n16091_ & ~new_n16422_;
  assign new_n16424_ = lo0234 & ~lo0505;
  assign new_n16425_ = ~new_n16118_ & ~new_n16424_;
  assign new_n16426_ = new_n16423_ & new_n16425_;
  assign new_n16427_ = new_n16411_ & new_n16416_;
  assign new_n16428_ = new_n16421_ & new_n16427_;
  assign new_n16429_ = new_n16426_ & new_n16428_;
  assign new_n16430_ = lo0240 & ~lo0542;
  assign new_n16431_ = ~new_n16229_ & ~new_n16430_;
  assign new_n16432_ = lo0244 & ~lo0541;
  assign new_n16433_ = ~new_n16226_ & ~new_n16432_;
  assign new_n16434_ = lo0242 & ~lo0539;
  assign new_n16435_ = ~new_n16220_ & ~new_n16434_;
  assign new_n16436_ = lo0245 & ~lo0503;
  assign new_n16437_ = ~new_n16112_ & ~new_n16436_;
  assign new_n16438_ = new_n16431_ & new_n16433_;
  assign new_n16439_ = new_n16435_ & new_n16438_;
  assign new_n16440_ = new_n16437_ & new_n16439_;
  assign new_n16441_ = lo0246 & lo0536;
  assign new_n16442_ = ~lo0246 & ~lo0536;
  assign new_n16443_ = ~new_n16441_ & ~new_n16442_;
  assign new_n16444_ = new_n14213_ & ~new_n16443_;
  assign new_n16445_ = lo0247 & ~lo0508;
  assign new_n16446_ = ~new_n16127_ & ~new_n16445_;
  assign new_n16447_ = new_n16444_ & new_n16446_;
  assign new_n16448_ = lo0241 & ~lo0506;
  assign new_n16449_ = ~new_n16121_ & ~new_n16448_;
  assign new_n16450_ = lo0248 & ~lo0537;
  assign new_n16451_ = ~new_n16214_ & ~new_n16450_;
  assign new_n16452_ = new_n16449_ & new_n16451_;
  assign new_n16453_ = lo0238 & ~lo0507;
  assign new_n16454_ = ~new_n16124_ & ~new_n16453_;
  assign new_n16455_ = lo0249 & ~lo0538;
  assign new_n16456_ = ~new_n16217_ & ~new_n16455_;
  assign new_n16457_ = new_n16454_ & new_n16456_;
  assign new_n16458_ = lo0234 & ~lo0557;
  assign new_n16459_ = ~new_n16274_ & ~new_n16458_;
  assign new_n16460_ = lo0235 & ~lo0533;
  assign new_n16461_ = ~new_n16202_ & ~new_n16460_;
  assign new_n16462_ = new_n16459_ & new_n16461_;
  assign new_n16463_ = new_n16447_ & new_n16452_;
  assign new_n16464_ = new_n16457_ & new_n16463_;
  assign new_n16465_ = new_n16462_ & new_n16464_;
  assign new_n16466_ = lo0240 & ~lo0535;
  assign new_n16467_ = ~new_n16208_ & ~new_n16466_;
  assign new_n16468_ = lo0245 & ~lo0509;
  assign new_n16469_ = ~new_n16130_ & ~new_n16468_;
  assign new_n16470_ = lo0242 & ~lo0504;
  assign new_n16471_ = ~new_n16115_ & ~new_n16470_;
  assign new_n16472_ = lo0244 & ~lo0558;
  assign new_n16473_ = ~new_n16277_ & ~new_n16472_;
  assign new_n16474_ = new_n16467_ & new_n16469_;
  assign new_n16475_ = new_n16471_ & new_n16474_;
  assign new_n16476_ = new_n16473_ & new_n16475_;
  assign new_n16477_ = lo0239 & ~lo0534;
  assign new_n16478_ = ~new_n16205_ & ~new_n16477_;
  assign new_n16479_ = new_n16476_ & new_n16478_;
  assign new_n16480_ = new_n16465_ & new_n16479_;
  assign new_n16481_ = new_n16429_ & new_n16440_;
  assign new_n16482_ = new_n16404_ & new_n16481_;
  assign new_n16483_ = ~new_n16480_ & ~new_n16482_;
  assign new_n16484_ = lo0239 & ~lo0550;
  assign new_n16485_ = ~new_n16253_ & ~new_n16484_;
  assign new_n16486_ = lo0246 & lo0563;
  assign new_n16487_ = ~lo0246 & ~lo0563;
  assign new_n16488_ = ~new_n16486_ & ~new_n16487_;
  assign new_n16489_ = new_n14285_ & ~new_n16488_;
  assign new_n16490_ = lo0247 & ~lo0552;
  assign new_n16491_ = ~new_n16259_ & ~new_n16490_;
  assign new_n16492_ = new_n16489_ & new_n16491_;
  assign new_n16493_ = lo0241 & ~lo0553;
  assign new_n16494_ = ~new_n16262_ & ~new_n16493_;
  assign new_n16495_ = lo0248 & ~lo0554;
  assign new_n16496_ = ~new_n16265_ & ~new_n16495_;
  assign new_n16497_ = new_n16494_ & new_n16496_;
  assign new_n16498_ = lo0238 & ~lo0577;
  assign new_n16499_ = ~new_n16340_ & ~new_n16498_;
  assign new_n16500_ = lo0249 & ~lo0555;
  assign new_n16501_ = ~new_n16268_ & ~new_n16500_;
  assign new_n16502_ = new_n16499_ & new_n16501_;
  assign new_n16503_ = lo0235 & ~lo0549;
  assign new_n16504_ = ~new_n16250_ & ~new_n16503_;
  assign new_n16505_ = lo0234 & ~lo0485;
  assign new_n16506_ = ~new_n16058_ & ~new_n16505_;
  assign new_n16507_ = new_n16504_ & new_n16506_;
  assign new_n16508_ = new_n16492_ & new_n16497_;
  assign new_n16509_ = new_n16502_ & new_n16508_;
  assign new_n16510_ = new_n16507_ & new_n16509_;
  assign new_n16511_ = lo0240 & ~lo0551;
  assign new_n16512_ = ~new_n16256_ & ~new_n16511_;
  assign new_n16513_ = lo0245 & ~lo0580;
  assign new_n16514_ = ~new_n16349_ & ~new_n16513_;
  assign new_n16515_ = lo0242 & ~lo0489;
  assign new_n16516_ = ~new_n16070_ & ~new_n16515_;
  assign new_n16517_ = lo0244 & ~lo0486;
  assign new_n16518_ = ~new_n16061_ & ~new_n16517_;
  assign new_n16519_ = new_n16512_ & new_n16514_;
  assign new_n16520_ = new_n16516_ & new_n16519_;
  assign new_n16521_ = new_n16518_ & new_n16520_;
  assign new_n16522_ = lo0248 & lo0548;
  assign new_n16523_ = ~lo0248 & ~lo0548;
  assign new_n16524_ = ~new_n16522_ & ~new_n16523_;
  assign new_n16525_ = new_n14306_ & ~new_n16524_;
  assign new_n16526_ = lo0241 & ~lo0490;
  assign new_n16527_ = ~new_n16073_ & ~new_n16526_;
  assign new_n16528_ = new_n16525_ & new_n16527_;
  assign new_n16529_ = lo0247 & ~lo0547;
  assign new_n16530_ = ~new_n16244_ & ~new_n16529_;
  assign new_n16531_ = lo0246 & ~lo0546;
  assign new_n16532_ = ~new_n16241_ & ~new_n16531_;
  assign new_n16533_ = new_n16530_ & new_n16532_;
  assign new_n16534_ = lo0238 & ~lo0491;
  assign new_n16535_ = ~new_n16076_ & ~new_n16534_;
  assign new_n16536_ = lo0234 & ~lo0544;
  assign new_n16537_ = ~new_n16235_ & ~new_n16536_;
  assign new_n16538_ = new_n16535_ & new_n16537_;
  assign new_n16539_ = lo0249 & ~lo0484;
  assign new_n16540_ = ~new_n16055_ & ~new_n16539_;
  assign new_n16541_ = lo0235 & ~lo0495;
  assign new_n16542_ = ~new_n16088_ & ~new_n16541_;
  assign new_n16543_ = new_n16540_ & new_n16542_;
  assign new_n16544_ = new_n16528_ & new_n16533_;
  assign new_n16545_ = new_n16538_ & new_n16544_;
  assign new_n16546_ = new_n16543_ & new_n16545_;
  assign new_n16547_ = lo0242 & ~lo0483;
  assign new_n16548_ = ~new_n16052_ & ~new_n16547_;
  assign new_n16549_ = lo0240 & ~lo0492;
  assign new_n16550_ = ~new_n16079_ & ~new_n16549_;
  assign new_n16551_ = lo0244 & ~lo0493;
  assign new_n16552_ = ~new_n16082_ & ~new_n16551_;
  assign new_n16553_ = lo0245 & ~lo0545;
  assign new_n16554_ = ~new_n16238_ & ~new_n16553_;
  assign new_n16555_ = new_n16548_ & new_n16550_;
  assign new_n16556_ = new_n16552_ & new_n16555_;
  assign new_n16557_ = new_n16554_ & new_n16556_;
  assign new_n16558_ = lo0239 & ~lo0494;
  assign new_n16559_ = ~new_n16085_ & ~new_n16558_;
  assign new_n16560_ = new_n16557_ & new_n16559_;
  assign new_n16561_ = new_n16546_ & new_n16560_;
  assign new_n16562_ = new_n16510_ & new_n16521_;
  assign new_n16563_ = new_n16485_ & new_n16562_;
  assign new_n16564_ = ~new_n16561_ & ~new_n16563_;
  assign new_n16565_ = new_n16483_ & new_n16564_;
  assign new_n16566_ = ~new_n4469_ & ~new_n16565_;
  assign new_n16567_ = lo0246 & lo0520;
  assign new_n16568_ = ~lo0246 & ~lo0520;
  assign new_n16569_ = ~new_n16567_ & ~new_n16568_;
  assign new_n16570_ = new_n14278_ & ~new_n16569_;
  assign new_n16571_ = lo0247 & ~lo0561;
  assign new_n16572_ = ~new_n16286_ & ~new_n16571_;
  assign new_n16573_ = new_n16570_ & new_n16572_;
  assign new_n16574_ = lo0241 & ~lo0574;
  assign new_n16575_ = ~new_n16331_ & ~new_n16574_;
  assign new_n16576_ = lo0248 & ~lo0521;
  assign new_n16577_ = ~new_n16166_ & ~new_n16576_;
  assign new_n16578_ = new_n16575_ & new_n16577_;
  assign new_n16579_ = lo0234 & ~lo0518;
  assign new_n16580_ = ~new_n16157_ & ~new_n16579_;
  assign new_n16581_ = lo0238 & ~lo0522;
  assign new_n16582_ = ~new_n16169_ & ~new_n16581_;
  assign new_n16583_ = new_n16580_ & new_n16582_;
  assign new_n16584_ = lo0249 & ~lo0578;
  assign new_n16585_ = ~new_n16343_ & ~new_n16584_;
  assign new_n16586_ = lo0235 & ~lo0581;
  assign new_n16587_ = ~new_n16352_ & ~new_n16586_;
  assign new_n16588_ = new_n16585_ & new_n16587_;
  assign new_n16589_ = new_n16573_ & new_n16578_;
  assign new_n16590_ = new_n16583_ & new_n16589_;
  assign new_n16591_ = new_n16588_ & new_n16590_;
  assign new_n16592_ = lo0245 & ~lo0584;
  assign new_n16593_ = ~new_n16358_ & ~new_n16592_;
  assign new_n16594_ = lo0240 & ~lo0582;
  assign new_n16595_ = ~new_n16355_ & ~new_n16594_;
  assign new_n16596_ = lo0244 & ~lo0585;
  assign new_n16597_ = ~new_n16361_ & ~new_n16596_;
  assign new_n16598_ = lo0242 & ~lo0586;
  assign new_n16599_ = ~new_n16364_ & ~new_n16598_;
  assign new_n16600_ = new_n16593_ & new_n16595_;
  assign new_n16601_ = new_n16597_ & new_n16600_;
  assign new_n16602_ = new_n16599_ & new_n16601_;
  assign new_n16603_ = new_n16591_ & new_n16602_;
  assign new_n16604_ = ~lo0239 & ~lo0519;
  assign new_n16605_ = lo0239 & lo0519;
  assign new_n16606_ = ~new_n16604_ & ~new_n16605_;
  assign new_n16607_ = lo0239 & ~lo0569;
  assign new_n16608_ = ~new_n16316_ & ~new_n16607_;
  assign new_n16609_ = lo0246 & lo0564;
  assign new_n16610_ = ~lo0246 & ~lo0564;
  assign new_n16611_ = ~new_n16609_ & ~new_n16610_;
  assign new_n16612_ = new_n14285_ & ~new_n16611_;
  assign new_n16613_ = lo0247 & ~lo0532;
  assign new_n16614_ = ~new_n16199_ & ~new_n16613_;
  assign new_n16615_ = new_n16612_ & new_n16614_;
  assign new_n16616_ = lo0248 & ~lo0565;
  assign new_n16617_ = ~new_n16298_ & ~new_n16616_;
  assign new_n16618_ = lo0241 & ~lo0562;
  assign new_n16619_ = ~new_n16289_ & ~new_n16618_;
  assign new_n16620_ = new_n16617_ & new_n16619_;
  assign new_n16621_ = lo0238 & ~lo0498;
  assign new_n16622_ = ~new_n16097_ & ~new_n16621_;
  assign new_n16623_ = lo0249 & ~lo0482;
  assign new_n16624_ = ~new_n16049_ & ~new_n16623_;
  assign new_n16625_ = new_n16622_ & new_n16624_;
  assign new_n16626_ = lo0234 & ~lo0570;
  assign new_n16627_ = ~new_n16319_ & ~new_n16626_;
  assign new_n16628_ = lo0235 & ~lo0531;
  assign new_n16629_ = ~new_n16196_ & ~new_n16628_;
  assign new_n16630_ = new_n16627_ & new_n16629_;
  assign new_n16631_ = new_n16615_ & new_n16620_;
  assign new_n16632_ = new_n16625_ & new_n16631_;
  assign new_n16633_ = new_n16630_ & new_n16632_;
  assign new_n16634_ = lo0240 & ~lo0560;
  assign new_n16635_ = ~new_n16283_ & ~new_n16634_;
  assign new_n16636_ = lo0245 & ~lo0568;
  assign new_n16637_ = ~new_n16313_ & ~new_n16636_;
  assign new_n16638_ = lo0242 & ~lo0556;
  assign new_n16639_ = ~new_n16271_ & ~new_n16638_;
  assign new_n16640_ = lo0244 & ~lo0566;
  assign new_n16641_ = ~new_n16301_ & ~new_n16640_;
  assign new_n16642_ = new_n16635_ & new_n16637_;
  assign new_n16643_ = new_n16639_ & new_n16642_;
  assign new_n16644_ = new_n16641_ & new_n16643_;
  assign new_n16645_ = lo0247 & lo0527;
  assign new_n16646_ = ~lo0247 & ~lo0527;
  assign new_n16647_ = ~new_n16645_ & ~new_n16646_;
  assign new_n16648_ = new_n14306_ & ~new_n16647_;
  assign new_n16649_ = lo0248 & ~lo0576;
  assign new_n16650_ = ~new_n16337_ & ~new_n16649_;
  assign new_n16651_ = new_n16648_ & new_n16650_;
  assign new_n16652_ = lo0246 & ~lo0526;
  assign new_n16653_ = ~new_n16181_ & ~new_n16652_;
  assign new_n16654_ = lo0241 & ~lo0571;
  assign new_n16655_ = ~new_n16322_ & ~new_n16654_;
  assign new_n16656_ = new_n16653_ & new_n16655_;
  assign new_n16657_ = lo0249 & ~lo0528;
  assign new_n16658_ = ~new_n16187_ & ~new_n16657_;
  assign new_n16659_ = lo0234 & ~lo0523;
  assign new_n16660_ = ~new_n16172_ & ~new_n16659_;
  assign new_n16661_ = new_n16658_ & new_n16660_;
  assign new_n16662_ = lo0235 & ~lo0575;
  assign new_n16663_ = ~new_n16334_ & ~new_n16662_;
  assign new_n16664_ = lo0238 & ~lo0529;
  assign new_n16665_ = ~new_n16190_ & ~new_n16664_;
  assign new_n16666_ = new_n16663_ & new_n16665_;
  assign new_n16667_ = new_n16651_ & new_n16656_;
  assign new_n16668_ = new_n16661_ & new_n16667_;
  assign new_n16669_ = new_n16666_ & new_n16668_;
  assign new_n16670_ = lo0240 & ~lo0530;
  assign new_n16671_ = ~new_n16193_ & ~new_n16670_;
  assign new_n16672_ = lo0245 & ~lo0525;
  assign new_n16673_ = ~new_n16178_ & ~new_n16672_;
  assign new_n16674_ = lo0242 & ~lo0573;
  assign new_n16675_ = ~new_n16328_ & ~new_n16674_;
  assign new_n16676_ = lo0244 & ~lo0572;
  assign new_n16677_ = ~new_n16325_ & ~new_n16676_;
  assign new_n16678_ = new_n16671_ & new_n16673_;
  assign new_n16679_ = new_n16675_ & new_n16678_;
  assign new_n16680_ = new_n16677_ & new_n16679_;
  assign new_n16681_ = lo0239 & ~lo0524;
  assign new_n16682_ = ~new_n16175_ & ~new_n16681_;
  assign new_n16683_ = new_n16680_ & new_n16682_;
  assign new_n16684_ = new_n16669_ & new_n16683_;
  assign new_n16685_ = new_n16633_ & new_n16644_;
  assign new_n16686_ = new_n16608_ & new_n16685_;
  assign new_n16687_ = ~new_n16684_ & ~new_n16686_;
  assign new_n16688_ = new_n16603_ & ~new_n16606_;
  assign new_n16689_ = new_n16687_ & ~new_n16688_;
  assign new_n16690_ = lo0247 & ~lo0516;
  assign new_n16691_ = ~new_n16151_ & ~new_n16690_;
  assign new_n16692_ = lo0248 & ~lo0481;
  assign new_n16693_ = ~new_n16046_ & ~new_n16692_;
  assign new_n16694_ = new_n16691_ & new_n16693_;
  assign new_n16695_ = lo0235 & ~lo0512;
  assign new_n16696_ = ~new_n16139_ & ~new_n16695_;
  assign new_n16697_ = lo0238 & ~lo0517;
  assign new_n16698_ = ~new_n16154_ & ~new_n16697_;
  assign new_n16699_ = new_n16696_ & new_n16698_;
  assign new_n16700_ = lo0234 & ~lo0511;
  assign new_n16701_ = ~new_n16136_ & ~new_n16700_;
  assign new_n16702_ = lo0249 & ~lo0579;
  assign new_n16703_ = ~new_n16346_ & ~new_n16702_;
  assign new_n16704_ = new_n16701_ & new_n16703_;
  assign new_n16705_ = new_n16694_ & new_n16699_;
  assign new_n16706_ = new_n16704_ & new_n16705_;
  assign new_n16707_ = lo0241 & lo0559;
  assign new_n16708_ = ~lo0241 & ~lo0559;
  assign new_n16709_ = ~new_n16707_ & ~new_n16708_;
  assign new_n16710_ = lo0246 & lo0487;
  assign new_n16711_ = ~lo0246 & ~lo0487;
  assign new_n16712_ = ~new_n16710_ & ~new_n16711_;
  assign new_n16713_ = ~new_n16709_ & ~new_n16712_;
  assign new_n16714_ = new_n14213_ & new_n16713_;
  assign new_n16715_ = new_n16706_ & new_n16714_;
  assign new_n16716_ = ~lo0239 & ~lo0488;
  assign new_n16717_ = lo0239 & lo0488;
  assign new_n16718_ = ~new_n16716_ & ~new_n16717_;
  assign new_n16719_ = lo0245 & ~lo0514;
  assign new_n16720_ = ~new_n16145_ & ~new_n16719_;
  assign new_n16721_ = lo0242 & ~lo0510;
  assign new_n16722_ = ~new_n16133_ & ~new_n16721_;
  assign new_n16723_ = new_n16720_ & new_n16722_;
  assign new_n16724_ = lo0240 & ~lo0515;
  assign new_n16725_ = ~new_n16148_ & ~new_n16724_;
  assign new_n16726_ = lo0244 & ~lo0513;
  assign new_n16727_ = ~new_n16142_ & ~new_n16726_;
  assign new_n16728_ = new_n16725_ & new_n16727_;
  assign new_n16729_ = new_n16715_ & ~new_n16718_;
  assign new_n16730_ = new_n16723_ & new_n16729_;
  assign new_n16731_ = new_n16728_ & new_n16730_;
  assign new_n16732_ = new_n16689_ & ~new_n16731_;
  assign new_n16733_ = new_n4460_ & ~new_n16732_;
  assign li0593 = new_n16566_ | new_n16733_;
  assign new_n16735_ = ~lo0594 & ~new_n15866_;
  assign new_n16736_ = ~new_n15867_ & ~new_n16735_;
  assign new_n16737_ = lo0806 & new_n16736_;
  assign new_n16738_ = lo0594 & ~lo0806;
  assign new_n16739_ = ~new_n16737_ & ~new_n16738_;
  assign li0594 = ~lo0332 & ~new_n16739_;
  assign new_n16741_ = lo0605 & new_n15860_;
  assign new_n16742_ = new_n15872_ & new_n16741_;
  assign new_n16743_ = ~lo0595 & ~new_n16742_;
  assign new_n16744_ = lo0595 & new_n16742_;
  assign new_n16745_ = ~new_n16743_ & ~new_n16744_;
  assign new_n16746_ = lo0806 & new_n16745_;
  assign new_n16747_ = lo0595 & ~lo0806;
  assign new_n16748_ = ~new_n16746_ & ~new_n16747_;
  assign li0595 = ~lo0332 & ~new_n16748_;
  assign new_n16750_ = new_n15895_ & new_n15897_;
  assign new_n16751_ = new_n15865_ & new_n16750_;
  assign new_n16752_ = ~lo0596 & ~new_n16751_;
  assign new_n16753_ = lo0596 & new_n16751_;
  assign new_n16754_ = ~new_n16752_ & ~new_n16753_;
  assign new_n16755_ = lo0806 & new_n16754_;
  assign new_n16756_ = lo0596 & ~lo0806;
  assign new_n16757_ = ~new_n16755_ & ~new_n16756_;
  assign li0596 = ~lo0332 & ~new_n16757_;
  assign new_n16759_ = lo0597 & new_n15867_;
  assign new_n16760_ = ~lo0597 & ~new_n15867_;
  assign new_n16761_ = ~new_n16759_ & ~new_n16760_;
  assign new_n16762_ = lo0806 & new_n16761_;
  assign new_n16763_ = lo0597 & ~lo0806;
  assign new_n16764_ = ~new_n16762_ & ~new_n16763_;
  assign li0597 = ~lo0332 & ~new_n16764_;
  assign li0882 = ~new_n3634_ | ~new_n4151_;
  assign new_n16767_ = lo0882 & ~li0882;
  assign new_n16768_ = lo0947 & new_n16767_;
  assign new_n16769_ = lo0598 & ~new_n16768_;
  assign new_n16770_ = lo0740 & ~lo0780;
  assign new_n16771_ = lo0603 & new_n16770_;
  assign new_n16772_ = new_n4453_ & new_n16771_;
  assign li0598 = new_n16769_ | new_n16772_;
  assign new_n16774_ = new_n15866_ & new_n15872_;
  assign new_n16775_ = new_n15885_ & new_n16774_;
  assign new_n16776_ = ~lo0599 & ~new_n16775_;
  assign new_n16777_ = lo0599 & new_n16775_;
  assign new_n16778_ = ~new_n16776_ & ~new_n16777_;
  assign new_n16779_ = lo0806 & new_n16778_;
  assign new_n16780_ = lo0599 & ~lo0806;
  assign new_n16781_ = ~new_n16779_ & ~new_n16780_;
  assign li0599 = ~lo0332 & ~new_n16781_;
  assign new_n16783_ = ~lo0600 & ~new_n15865_;
  assign new_n16784_ = ~new_n15866_ & ~new_n16783_;
  assign new_n16785_ = lo0806 & new_n16784_;
  assign new_n16786_ = lo0600 & ~lo0806;
  assign new_n16787_ = ~new_n16785_ & ~new_n16786_;
  assign li0600 = ~lo0332 & ~new_n16787_;
  assign new_n16789_ = lo0601 & ~lo0806;
  assign new_n16790_ = lo0601 & ~lo0605;
  assign new_n16791_ = ~lo0601 & lo0605;
  assign new_n16792_ = ~new_n16790_ & ~new_n16791_;
  assign new_n16793_ = lo0806 & ~new_n16792_;
  assign new_n16794_ = ~new_n16789_ & ~new_n16793_;
  assign li0601 = ~lo0332 & ~new_n16794_;
  assign new_n16796_ = lo0230 & lo0602;
  assign new_n16797_ = ~lo0602 & new_n13786_;
  assign li0602 = new_n16796_ | new_n16797_;
  assign new_n16799_ = lo0871 & lo0966;
  assign new_n16800_ = ~lo0980 & lo1055;
  assign new_n16801_ = ~lo1032 & new_n16800_;
  assign new_n16802_ = lo0832 & new_n16801_;
  assign new_n16803_ = ~lo1054 & new_n16802_;
  assign li0740 = ~lo0952 & new_n16803_;
  assign new_n16805_ = pi011 & li0740;
  assign new_n16806_ = lo0603 & ~li0740;
  assign new_n16807_ = ~new_n16805_ & ~new_n16806_;
  assign new_n16808_ = ~lo0966 & ~new_n16807_;
  assign new_n16809_ = lo0872 & lo0966;
  assign new_n16810_ = ~new_n16799_ & ~new_n16808_;
  assign li0603 = new_n16809_ | ~new_n16810_;
  assign new_n16812_ = ~lo0661 & new_n4465_;
  assign new_n16813_ = lo0823 & new_n16812_;
  assign new_n16814_ = lo0779 & new_n16813_;
  assign new_n16815_ = ~lo0299 & lo0983;
  assign new_n16816_ = lo0907 & new_n16815_;
  assign new_n16817_ = ~new_n16813_ & ~new_n16816_;
  assign new_n16818_ = lo0604 & new_n16817_;
  assign li0604 = new_n16814_ | new_n16818_;
  assign new_n16820_ = ~lo0605 & ~lo0806;
  assign new_n16821_ = lo0605 & lo0806;
  assign new_n16822_ = ~new_n16820_ & ~new_n16821_;
  assign li0605 = ~lo0332 & new_n16822_;
  assign new_n16824_ = pi015 & ~li0740;
  assign new_n16825_ = ~pi015 & lo0606;
  assign new_n16826_ = ~new_n16824_ & ~new_n16825_;
  assign new_n16827_ = lo0966 & ~new_n16826_;
  assign new_n16828_ = lo0837 & new_n16826_;
  assign li0606 = new_n16827_ | new_n16828_;
  assign new_n16830_ = lo0607 & ~li0740;
  assign new_n16831_ = pi018 & li0740;
  assign new_n16832_ = ~new_n16830_ & ~new_n16831_;
  assign li0607 = ~lo0966 & ~new_n16832_;
  assign new_n16834_ = lo0608 & ~li0740;
  assign new_n16835_ = pi027 & li0740;
  assign new_n16836_ = ~new_n16834_ & ~new_n16835_;
  assign li0608 = ~lo0966 & ~new_n16836_;
  assign new_n16838_ = lo0609 & ~li0740;
  assign new_n16839_ = pi029 & li0740;
  assign new_n16840_ = ~new_n16838_ & ~new_n16839_;
  assign li0609 = ~lo0966 & ~new_n16840_;
  assign new_n16842_ = lo0610 & ~li0740;
  assign new_n16843_ = pi024 & li0740;
  assign new_n16844_ = ~new_n16842_ & ~new_n16843_;
  assign li0610 = ~lo0966 & ~new_n16844_;
  assign new_n16846_ = lo0611 & ~li0740;
  assign new_n16847_ = pi025 & li0740;
  assign new_n16848_ = ~new_n16846_ & ~new_n16847_;
  assign li0611 = ~lo0966 & ~new_n16848_;
  assign new_n16850_ = lo0612 & ~li0740;
  assign new_n16851_ = pi022 & li0740;
  assign new_n16852_ = ~new_n16850_ & ~new_n16851_;
  assign li0612 = ~lo0966 & ~new_n16852_;
  assign new_n16854_ = lo0613 & ~li0740;
  assign new_n16855_ = pi026 & li0740;
  assign new_n16856_ = ~new_n16854_ & ~new_n16855_;
  assign li0613 = ~lo0966 & ~new_n16856_;
  assign new_n16858_ = pi013 & li0740;
  assign new_n16859_ = lo0614 & ~li0740;
  assign new_n16860_ = ~new_n16858_ & ~new_n16859_;
  assign new_n16861_ = ~lo0966 & ~new_n16860_;
  assign li0614 = new_n16799_ | new_n16861_;
  assign new_n16863_ = lo0907 & new_n16767_;
  assign new_n16864_ = ~lo0779 & lo0797;
  assign new_n16865_ = lo0680 & new_n16864_;
  assign new_n16866_ = new_n16812_ & new_n16865_;
  assign new_n16867_ = lo0615 & ~new_n16863_;
  assign li0615 = new_n16866_ | new_n16867_;
  assign new_n16869_ = pi012 & li0740;
  assign new_n16870_ = lo0616 & ~li0740;
  assign new_n16871_ = ~new_n16869_ & ~new_n16870_;
  assign new_n16872_ = ~lo0966 & ~new_n16871_;
  assign li0616 = new_n16809_ | new_n16872_;
  assign new_n16874_ = pi016 & ~li0740;
  assign new_n16875_ = ~pi016 & lo0617;
  assign new_n16876_ = ~new_n16874_ & ~new_n16875_;
  assign new_n16877_ = lo0966 & ~new_n16876_;
  assign new_n16878_ = lo0850 & new_n16876_;
  assign li0617 = new_n16877_ | new_n16878_;
  assign new_n16880_ = lo0618 & ~li0740;
  assign new_n16881_ = pi028 & li0740;
  assign new_n16882_ = ~new_n16880_ & ~new_n16881_;
  assign li0618 = ~lo0966 & ~new_n16882_;
  assign new_n16884_ = lo0619 & ~li0740;
  assign new_n16885_ = pi033 & li0740;
  assign new_n16886_ = ~new_n16884_ & ~new_n16885_;
  assign li0619 = ~lo0966 & ~new_n16886_;
  assign new_n16888_ = lo0620 & ~li0740;
  assign new_n16889_ = pi023 & li0740;
  assign new_n16890_ = ~new_n16888_ & ~new_n16889_;
  assign li0620 = ~lo0966 & ~new_n16890_;
  assign new_n16892_ = lo0621 & ~li0740;
  assign new_n16893_ = pi019 & li0740;
  assign new_n16894_ = ~new_n16892_ & ~new_n16893_;
  assign li0621 = ~lo0966 & ~new_n16894_;
  assign new_n16896_ = lo0622 & ~li0740;
  assign new_n16897_ = pi020 & li0740;
  assign new_n16898_ = ~new_n16896_ & ~new_n16897_;
  assign li0622 = ~lo0966 & ~new_n16898_;
  assign new_n16900_ = lo0623 & ~li0740;
  assign new_n16901_ = pi017 & li0740;
  assign new_n16902_ = ~new_n16900_ & ~new_n16901_;
  assign li0623 = ~lo0966 & ~new_n16902_;
  assign new_n16904_ = lo0831 & new_n4453_;
  assign new_n16905_ = lo0780 & new_n16904_;
  assign new_n16906_ = lo0947 & new_n16815_;
  assign new_n16907_ = ~new_n16904_ & ~new_n16906_;
  assign new_n16908_ = lo0624 & new_n16907_;
  assign li0624 = new_n16905_ | new_n16908_;
  assign new_n16910_ = lo0973 & lo1048;
  assign new_n16911_ = ~lo1082 & new_n16910_;
  assign new_n16912_ = lo0832 & new_n16911_;
  assign new_n16913_ = ~lo1060 & new_n16912_;
  assign li0797 = ~lo0953 & new_n16913_;
  assign new_n16915_ = lo0625 & ~li0797;
  assign new_n16916_ = pi027 & li0797;
  assign new_n16917_ = ~new_n16915_ & ~new_n16916_;
  assign li0625 = ~lo0962 & ~new_n16917_;
  assign new_n16919_ = lo0626 & ~li0740;
  assign new_n16920_ = pi032 & li0740;
  assign new_n16921_ = ~new_n16919_ & ~new_n16920_;
  assign li0626 = ~lo0966 & ~new_n16921_;
  assign new_n16923_ = lo0627 & ~li0797;
  assign new_n16924_ = pi028 & li0797;
  assign new_n16925_ = ~new_n16923_ & ~new_n16924_;
  assign li0627 = ~lo0962 & ~new_n16925_;
  assign new_n16927_ = lo0628 & ~li0797;
  assign new_n16928_ = pi030 & li0797;
  assign new_n16929_ = ~new_n16927_ & ~new_n16928_;
  assign li0628 = ~lo0962 & ~new_n16929_;
  assign new_n16931_ = lo0629 & ~li0740;
  assign new_n16932_ = pi030 & li0740;
  assign new_n16933_ = ~new_n16931_ & ~new_n16932_;
  assign li0629 = ~lo0966 & ~new_n16933_;
  assign new_n16935_ = lo0630 & ~li0740;
  assign new_n16936_ = pi031 & li0740;
  assign new_n16937_ = ~new_n16935_ & ~new_n16936_;
  assign li0630 = ~lo0966 & ~new_n16937_;
  assign new_n16939_ = lo0631 & ~li0797;
  assign new_n16940_ = pi024 & li0797;
  assign new_n16941_ = ~new_n16939_ & ~new_n16940_;
  assign li0631 = ~lo0962 & ~new_n16941_;
  assign new_n16943_ = lo0632 & ~li0797;
  assign new_n16944_ = pi026 & li0797;
  assign new_n16945_ = ~new_n16943_ & ~new_n16944_;
  assign li0632 = ~lo0962 & ~new_n16945_;
  assign new_n16947_ = lo0633 & ~li0740;
  assign new_n16948_ = pi021 & li0740;
  assign new_n16949_ = ~new_n16947_ & ~new_n16948_;
  assign li0633 = ~lo0966 & ~new_n16949_;
  assign new_n16951_ = lo0634 & ~li0797;
  assign new_n16952_ = pi021 & li0797;
  assign new_n16953_ = ~new_n16951_ & ~new_n16952_;
  assign li0634 = ~lo0962 & ~new_n16953_;
  assign new_n16955_ = lo0635 & ~li0797;
  assign new_n16956_ = pi023 & li0797;
  assign new_n16957_ = ~new_n16955_ & ~new_n16956_;
  assign li0635 = ~lo0962 & ~new_n16957_;
  assign new_n16959_ = lo0636 & ~li0740;
  assign new_n16960_ = pi038 & li0740;
  assign new_n16961_ = ~new_n16959_ & ~new_n16960_;
  assign li0636 = ~lo0966 & ~new_n16961_;
  assign new_n16963_ = lo0637 & ~li0797;
  assign new_n16964_ = pi016 & li0797;
  assign new_n16965_ = ~new_n16963_ & ~new_n16964_;
  assign li0637 = ~lo0962 & ~new_n16965_;
  assign new_n16967_ = lo0638 & ~li0797;
  assign new_n16968_ = pi018 & li0797;
  assign new_n16969_ = ~new_n16967_ & ~new_n16968_;
  assign li0638 = ~lo0962 & ~new_n16969_;
  assign new_n16971_ = lo0639 & ~li0797;
  assign new_n16972_ = pi020 & li0797;
  assign new_n16973_ = ~new_n16971_ & ~new_n16972_;
  assign li0639 = ~lo0962 & ~new_n16973_;
  assign new_n16975_ = lo0640 & ~li0740;
  assign new_n16976_ = pi039 & li0740;
  assign new_n16977_ = ~new_n16975_ & ~new_n16976_;
  assign li0640 = ~lo0966 & ~new_n16977_;
  assign new_n16979_ = lo0641 & ~li0797;
  assign new_n16980_ = pi032 & li0797;
  assign new_n16981_ = ~new_n16979_ & ~new_n16980_;
  assign li0641 = ~lo0962 & ~new_n16981_;
  assign new_n16983_ = lo0642 & ~li0740;
  assign new_n16984_ = pi014 & li0740;
  assign new_n16985_ = ~new_n16983_ & ~new_n16984_;
  assign li0642 = ~lo0966 & ~new_n16985_;
  assign new_n16987_ = lo0643 & ~li0797;
  assign new_n16988_ = pi015 & li0797;
  assign new_n16989_ = ~new_n16987_ & ~new_n16988_;
  assign li0643 = ~lo0962 & ~new_n16989_;
  assign new_n16991_ = lo0644 & ~li0740;
  assign new_n16992_ = pi034 & li0740;
  assign new_n16993_ = ~new_n16991_ & ~new_n16992_;
  assign li0644 = ~lo0966 & ~new_n16993_;
  assign new_n16995_ = lo0645 & ~li0740;
  assign new_n16996_ = pi036 & li0740;
  assign new_n16997_ = ~new_n16995_ & ~new_n16996_;
  assign li0645 = ~lo0966 & ~new_n16997_;
  assign new_n16999_ = lo0646 & ~li0797;
  assign new_n17000_ = pi025 & li0797;
  assign new_n17001_ = ~new_n16999_ & ~new_n17000_;
  assign li0646 = ~lo0962 & ~new_n17001_;
  assign new_n17003_ = lo0647 & ~li0797;
  assign new_n17004_ = pi031 & li0797;
  assign new_n17005_ = ~new_n17003_ & ~new_n17004_;
  assign li0647 = ~lo0962 & ~new_n17005_;
  assign new_n17007_ = lo0648 & ~li0797;
  assign new_n17008_ = pi033 & li0797;
  assign new_n17009_ = ~new_n17007_ & ~new_n17008_;
  assign li0648 = ~lo0962 & ~new_n17009_;
  assign new_n17011_ = lo0649 & ~li0797;
  assign new_n17012_ = pi037 & li0797;
  assign new_n17013_ = ~new_n17011_ & ~new_n17012_;
  assign li0649 = ~lo0962 & ~new_n17013_;
  assign new_n17015_ = lo0650 & ~li0797;
  assign new_n17016_ = pi038 & li0797;
  assign new_n17017_ = ~new_n17015_ & ~new_n17016_;
  assign li0650 = ~lo0962 & ~new_n17017_;
  assign new_n17019_ = lo0651 & ~li0740;
  assign new_n17020_ = pi041 & li0740;
  assign new_n17021_ = ~new_n17019_ & ~new_n17020_;
  assign li0651 = ~lo0966 & ~new_n17021_;
  assign new_n17023_ = lo0652 & ~li0740;
  assign new_n17024_ = pi042 & li0740;
  assign new_n17025_ = ~new_n17023_ & ~new_n17024_;
  assign li0652 = ~lo0966 & ~new_n17025_;
  assign new_n17027_ = lo0653 & ~li0740;
  assign new_n17028_ = pi040 & li0740;
  assign new_n17029_ = ~new_n17027_ & ~new_n17028_;
  assign li0653 = ~lo0966 & ~new_n17029_;
  assign new_n17031_ = lo0654 & ~li0797;
  assign new_n17032_ = pi041 & li0797;
  assign new_n17033_ = ~new_n17031_ & ~new_n17032_;
  assign li0654 = ~lo0962 & ~new_n17033_;
  assign new_n17035_ = lo0655 & ~li0797;
  assign new_n17036_ = pi035 & li0797;
  assign new_n17037_ = ~new_n17035_ & ~new_n17036_;
  assign li0655 = ~lo0962 & ~new_n17037_;
  assign new_n17039_ = lo0656 & ~li0740;
  assign new_n17040_ = pi037 & li0740;
  assign new_n17041_ = ~new_n17039_ & ~new_n17040_;
  assign li0656 = ~lo0966 & ~new_n17041_;
  assign new_n17043_ = lo0657 & ~li0797;
  assign new_n17044_ = pi042 & li0797;
  assign new_n17045_ = ~new_n17043_ & ~new_n17044_;
  assign li0657 = ~lo0962 & ~new_n17045_;
  assign new_n17047_ = lo0658 & ~li0740;
  assign new_n17048_ = pi035 & li0740;
  assign new_n17049_ = ~new_n17047_ & ~new_n17048_;
  assign li0658 = ~lo0966 & ~new_n17049_;
  assign new_n17051_ = lo0278 & lo0279;
  assign new_n17052_ = lo0266 & new_n17051_;
  assign new_n17053_ = lo0280 & new_n17052_;
  assign new_n17054_ = lo0269 & new_n17053_;
  assign new_n17055_ = lo0282 & new_n17054_;
  assign new_n17056_ = lo0281 & new_n17055_;
  assign new_n17057_ = lo0264 & lo0277;
  assign new_n17058_ = new_n17056_ & new_n17057_;
  assign new_n17059_ = lo0265 & new_n17058_;
  assign new_n17060_ = lo0270 & new_n17059_;
  assign new_n17061_ = lo0274 & ~new_n17060_;
  assign new_n17062_ = ~lo0274 & new_n17060_;
  assign li0659 = new_n17061_ | new_n17062_;
  assign new_n17064_ = lo0660 & ~li0797;
  assign new_n17065_ = pi029 & li0797;
  assign new_n17066_ = ~new_n17064_ & ~new_n17065_;
  assign li0660 = ~lo0962 & ~new_n17066_;
  assign new_n17068_ = lo0661 & ~li0797;
  assign new_n17069_ = pi012 & li0797;
  assign new_n17070_ = ~new_n17068_ & ~new_n17069_;
  assign li0661 = ~lo0962 & ~new_n17070_;
  assign new_n17072_ = lo0662 & ~li0797;
  assign new_n17073_ = pi013 & li0797;
  assign new_n17074_ = ~new_n17072_ & ~new_n17073_;
  assign li0662 = ~lo0962 & ~new_n17074_;
  assign new_n17076_ = ~pi048 & ~pi049;
  assign new_n17077_ = ~pi046 & new_n17076_;
  assign new_n17078_ = pi047 & new_n17077_;
  assign new_n17079_ = pi045 & new_n17078_;
  assign new_n17080_ = ~pi045 & new_n17078_;
  assign new_n17081_ = lo0766 & new_n17079_;
  assign new_n17082_ = lo0633 & new_n17080_;
  assign new_n17083_ = ~new_n17081_ & ~new_n17082_;
  assign new_n17084_ = pi046 & new_n17076_;
  assign new_n17085_ = pi047 & new_n17084_;
  assign new_n17086_ = pi045 & new_n17085_;
  assign new_n17087_ = ~pi045 & new_n17085_;
  assign new_n17088_ = lo0700 & new_n17086_;
  assign new_n17089_ = lo0634 & new_n17087_;
  assign new_n17090_ = ~new_n17088_ & ~new_n17089_;
  assign new_n17091_ = ~pi046 & ~pi047;
  assign new_n17092_ = new_n17076_ & new_n17091_;
  assign new_n17093_ = pi045 & new_n17092_;
  assign new_n17094_ = lo0855 & new_n17093_;
  assign new_n17095_ = ~pi045 & new_n17076_;
  assign new_n17096_ = pi046 & ~pi047;
  assign new_n17097_ = new_n17095_ & new_n17096_;
  assign new_n17098_ = ~pi045 & new_n17092_;
  assign new_n17099_ = lo0784 & new_n17097_;
  assign new_n17100_ = lo0815 & new_n17098_;
  assign new_n17101_ = ~new_n17099_ & ~new_n17100_;
  assign new_n17102_ = new_n17083_ & new_n17090_;
  assign new_n17103_ = ~new_n17094_ & new_n17102_;
  assign new_n17104_ = new_n17101_ & new_n17103_;
  assign new_n17105_ = ~new_n14878_ & ~new_n14883_;
  assign new_n17106_ = lo0257 & ~new_n17105_;
  assign new_n17107_ = lo0199 & lo1059;
  assign new_n17108_ = ~new_n17106_ & ~new_n17107_;
  assign new_n17109_ = ~lo0223 & ~lo0224;
  assign new_n17110_ = lo0222 & new_n17109_;
  assign new_n17111_ = ~lo0222 & ~lo0223;
  assign new_n17112_ = ~lo0224 & new_n17111_;
  assign new_n17113_ = ~new_n17110_ & ~new_n17112_;
  assign new_n17114_ = ~new_n5022_ & ~new_n17113_;
  assign new_n17115_ = ~new_n17108_ & new_n17113_;
  assign new_n17116_ = ~new_n17114_ & ~new_n17115_;
  assign new_n17117_ = new_n5051_ & ~new_n17104_;
  assign new_n17118_ = new_n17104_ & ~new_n17116_;
  assign li0663 = new_n17117_ | new_n17118_;
  assign new_n17120_ = lo0772 & new_n17079_;
  assign new_n17121_ = lo0614 & new_n17080_;
  assign new_n17122_ = ~new_n17120_ & ~new_n17121_;
  assign new_n17123_ = lo0727 & new_n17086_;
  assign new_n17124_ = lo0662 & new_n17087_;
  assign new_n17125_ = ~new_n17123_ & ~new_n17124_;
  assign new_n17126_ = lo0811 & new_n17098_;
  assign new_n17127_ = lo0785 & new_n17097_;
  assign new_n17128_ = lo0872 & new_n17093_;
  assign new_n17129_ = ~new_n17127_ & ~new_n17128_;
  assign new_n17130_ = new_n17122_ & new_n17125_;
  assign new_n17131_ = ~new_n17126_ & new_n17130_;
  assign new_n17132_ = new_n17129_ & new_n17131_;
  assign new_n17133_ = lo0292 & ~new_n17105_;
  assign new_n17134_ = lo0199 & lo1078;
  assign new_n17135_ = ~new_n17133_ & ~new_n17134_;
  assign new_n17136_ = ~new_n4721_ & ~new_n17113_;
  assign new_n17137_ = new_n17113_ & ~new_n17135_;
  assign new_n17138_ = ~new_n17136_ & ~new_n17137_;
  assign new_n17139_ = new_n5051_ & ~new_n17132_;
  assign new_n17140_ = new_n17132_ & ~new_n17138_;
  assign li0664 = new_n17139_ | new_n17140_;
  assign new_n17142_ = lo0665 & ~li0797;
  assign new_n17143_ = pi019 & li0797;
  assign new_n17144_ = ~new_n17142_ & ~new_n17143_;
  assign li0665 = ~lo0962 & ~new_n17144_;
  assign new_n17146_ = lo0764 & new_n17079_;
  assign new_n17147_ = lo0607 & new_n17080_;
  assign new_n17148_ = ~new_n17146_ & ~new_n17147_;
  assign new_n17149_ = lo0691 & new_n17086_;
  assign new_n17150_ = lo0638 & new_n17087_;
  assign new_n17151_ = ~new_n17149_ & ~new_n17150_;
  assign new_n17152_ = lo0873 & new_n17093_;
  assign new_n17153_ = lo0790 & new_n17097_;
  assign new_n17154_ = lo0799 & new_n17098_;
  assign new_n17155_ = ~new_n17153_ & ~new_n17154_;
  assign new_n17156_ = new_n17148_ & new_n17151_;
  assign new_n17157_ = ~new_n17152_ & new_n17156_;
  assign new_n17158_ = new_n17155_ & new_n17157_;
  assign new_n17159_ = lo0297 & ~new_n17105_;
  assign new_n17160_ = lo0199 & lo1038;
  assign new_n17161_ = ~new_n17159_ & ~new_n17160_;
  assign new_n17162_ = ~new_n4704_ & ~new_n17113_;
  assign new_n17163_ = new_n17113_ & ~new_n17161_;
  assign new_n17164_ = ~new_n17162_ & ~new_n17163_;
  assign new_n17165_ = new_n5051_ & ~new_n17158_;
  assign new_n17166_ = new_n17158_ & ~new_n17164_;
  assign li0666 = new_n17165_ | new_n17166_;
  assign new_n17168_ = lo0792 & new_n17097_;
  assign new_n17169_ = lo0871 & new_n17093_;
  assign new_n17170_ = ~new_n17168_ & ~new_n17169_;
  assign new_n17171_ = lo0809 & new_n17098_;
  assign new_n17172_ = lo0699 & new_n17086_;
  assign new_n17173_ = lo0681 & new_n17087_;
  assign new_n17174_ = ~new_n17172_ & ~new_n17173_;
  assign new_n17175_ = lo0763 & new_n17079_;
  assign new_n17176_ = lo0642 & new_n17080_;
  assign new_n17177_ = ~new_n17175_ & ~new_n17176_;
  assign new_n17178_ = new_n17170_ & ~new_n17171_;
  assign new_n17179_ = new_n17174_ & new_n17178_;
  assign new_n17180_ = new_n17177_ & new_n17179_;
  assign new_n17181_ = lo0294 & ~new_n17105_;
  assign new_n17182_ = lo0199 & lo1066;
  assign new_n17183_ = ~new_n17181_ & ~new_n17182_;
  assign new_n17184_ = ~new_n4741_ & ~new_n17113_;
  assign new_n17185_ = new_n17113_ & ~new_n17183_;
  assign new_n17186_ = ~new_n17184_ & ~new_n17185_;
  assign new_n17187_ = new_n5051_ & ~new_n17180_;
  assign new_n17188_ = new_n17180_ & ~new_n17186_;
  assign li0667 = new_n17187_ | new_n17188_;
  assign new_n17190_ = lo0759 & new_n17079_;
  assign new_n17191_ = lo0603 & new_n17080_;
  assign new_n17192_ = ~new_n17190_ & ~new_n17191_;
  assign new_n17193_ = lo0696 & new_n17086_;
  assign new_n17194_ = lo0680 & new_n17087_;
  assign new_n17195_ = ~new_n17193_ & ~new_n17194_;
  assign new_n17196_ = lo0837 & new_n17093_;
  assign new_n17197_ = lo0778 & new_n17097_;
  assign new_n17198_ = lo0981 & new_n17098_;
  assign new_n17199_ = ~new_n17197_ & ~new_n17198_;
  assign new_n17200_ = new_n17192_ & new_n17195_;
  assign new_n17201_ = ~new_n17196_ & new_n17200_;
  assign new_n17202_ = new_n17199_ & new_n17201_;
  assign new_n17203_ = lo0291 & ~new_n17105_;
  assign new_n17204_ = lo0199 & lo1043;
  assign new_n17205_ = ~new_n17203_ & ~new_n17204_;
  assign new_n17206_ = ~new_n4711_ & ~new_n17113_;
  assign new_n17207_ = new_n17113_ & ~new_n17205_;
  assign new_n17208_ = ~new_n17206_ & ~new_n17207_;
  assign new_n17209_ = new_n5051_ & ~new_n17202_;
  assign new_n17210_ = new_n17202_ & ~new_n17208_;
  assign li0668 = new_n17209_ | new_n17210_;
  assign new_n17212_ = lo0669 & ~li0797;
  assign new_n17213_ = pi036 & li0797;
  assign new_n17214_ = ~new_n17212_ & ~new_n17213_;
  assign li0669 = ~lo0962 & ~new_n17214_;
  assign new_n17216_ = lo0723 & new_n17086_;
  assign new_n17217_ = lo0695 & new_n17087_;
  assign new_n17218_ = ~new_n17216_ & ~new_n17217_;
  assign new_n17219_ = lo0745 & new_n17079_;
  assign new_n17220_ = lo0612 & new_n17080_;
  assign new_n17221_ = lo0852 & new_n17093_;
  assign new_n17222_ = ~new_n17220_ & ~new_n17221_;
  assign new_n17223_ = new_n17218_ & ~new_n17219_;
  assign new_n17224_ = new_n17222_ & new_n17223_;
  assign new_n17225_ = lo0258 & ~new_n17105_;
  assign new_n17226_ = lo0199 & lo1056;
  assign new_n17227_ = ~new_n17225_ & ~new_n17226_;
  assign new_n17228_ = ~new_n4968_ & ~new_n17113_;
  assign new_n17229_ = new_n17113_ & ~new_n17227_;
  assign new_n17230_ = ~new_n17228_ & ~new_n17229_;
  assign new_n17231_ = new_n5051_ & ~new_n17224_;
  assign new_n17232_ = new_n17224_ & ~new_n17230_;
  assign li0670 = new_n17231_ | new_n17232_;
  assign new_n17234_ = lo0724 & new_n17086_;
  assign new_n17235_ = lo0646 & new_n17087_;
  assign new_n17236_ = ~new_n17234_ & ~new_n17235_;
  assign new_n17237_ = lo0741 & new_n17079_;
  assign new_n17238_ = lo0611 & new_n17080_;
  assign new_n17239_ = lo0865 & new_n17093_;
  assign new_n17240_ = ~new_n17238_ & ~new_n17239_;
  assign new_n17241_ = new_n17236_ & ~new_n17237_;
  assign new_n17242_ = new_n17240_ & new_n17241_;
  assign new_n17243_ = lo0261 & ~new_n17105_;
  assign new_n17244_ = lo0199 & lo1034;
  assign new_n17245_ = ~new_n17243_ & ~new_n17244_;
  assign new_n17246_ = ~new_n4992_ & ~new_n17113_;
  assign new_n17247_ = new_n17113_ & ~new_n17245_;
  assign new_n17248_ = ~new_n17246_ & ~new_n17247_;
  assign new_n17249_ = new_n5051_ & ~new_n17242_;
  assign new_n17250_ = new_n17242_ & ~new_n17248_;
  assign li0671 = new_n17249_ | new_n17250_;
  assign new_n17252_ = lo0781 & new_n17097_;
  assign new_n17253_ = lo0850 & new_n17093_;
  assign new_n17254_ = ~new_n17252_ & ~new_n17253_;
  assign new_n17255_ = lo0808 & new_n17098_;
  assign new_n17256_ = lo0758 & new_n17079_;
  assign new_n17257_ = lo0616 & new_n17080_;
  assign new_n17258_ = ~new_n17256_ & ~new_n17257_;
  assign new_n17259_ = lo0736 & new_n17086_;
  assign new_n17260_ = lo0661 & new_n17087_;
  assign new_n17261_ = ~new_n17259_ & ~new_n17260_;
  assign new_n17262_ = new_n17254_ & ~new_n17255_;
  assign new_n17263_ = new_n17258_ & new_n17262_;
  assign new_n17264_ = new_n17261_ & new_n17263_;
  assign new_n17265_ = lo0290 & ~new_n17105_;
  assign new_n17266_ = lo0199 & lo1042;
  assign new_n17267_ = ~new_n17265_ & ~new_n17266_;
  assign new_n17268_ = ~new_n4758_ & ~new_n17113_;
  assign new_n17269_ = new_n17113_ & ~new_n17267_;
  assign new_n17270_ = ~new_n17268_ & ~new_n17269_;
  assign new_n17271_ = new_n5051_ & ~new_n17264_;
  assign new_n17272_ = new_n17264_ & ~new_n17270_;
  assign li0672 = new_n17271_ | new_n17272_;
  assign new_n17274_ = lo0788 & new_n17097_;
  assign new_n17275_ = lo0866 & new_n17093_;
  assign new_n17276_ = ~new_n17274_ & ~new_n17275_;
  assign new_n17277_ = lo0814 & new_n17098_;
  assign new_n17278_ = lo0706 & new_n17086_;
  assign new_n17279_ = lo0637 & new_n17087_;
  assign new_n17280_ = ~new_n17278_ & ~new_n17279_;
  assign new_n17281_ = lo0749 & new_n17079_;
  assign new_n17282_ = lo0617 & new_n17080_;
  assign new_n17283_ = ~new_n17281_ & ~new_n17282_;
  assign new_n17284_ = new_n17276_ & ~new_n17277_;
  assign new_n17285_ = new_n17280_ & new_n17284_;
  assign new_n17286_ = new_n17283_ & new_n17285_;
  assign new_n17287_ = lo0295 & ~new_n17105_;
  assign new_n17288_ = lo0199 & lo1047;
  assign new_n17289_ = ~new_n17287_ & ~new_n17288_;
  assign new_n17290_ = ~new_n4748_ & ~new_n17113_;
  assign new_n17291_ = new_n17113_ & ~new_n17289_;
  assign new_n17292_ = ~new_n17290_ & ~new_n17291_;
  assign new_n17293_ = new_n5051_ & ~new_n17286_;
  assign new_n17294_ = new_n17286_ & ~new_n17292_;
  assign li0673 = new_n17293_ | new_n17294_;
  assign new_n17296_ = lo0783 & new_n17097_;
  assign new_n17297_ = lo0859 & new_n17093_;
  assign new_n17298_ = ~new_n17296_ & ~new_n17297_;
  assign new_n17299_ = lo0804 & new_n17098_;
  assign new_n17300_ = lo0743 & new_n17079_;
  assign new_n17301_ = lo0622 & new_n17080_;
  assign new_n17302_ = ~new_n17300_ & ~new_n17301_;
  assign new_n17303_ = lo0735 & new_n17086_;
  assign new_n17304_ = lo0639 & new_n17087_;
  assign new_n17305_ = ~new_n17303_ & ~new_n17304_;
  assign new_n17306_ = new_n17298_ & ~new_n17299_;
  assign new_n17307_ = new_n17302_ & new_n17306_;
  assign new_n17308_ = new_n17305_ & new_n17307_;
  assign new_n17309_ = lo0256 & ~new_n17105_;
  assign new_n17310_ = lo0199 & lo1064;
  assign new_n17311_ = ~new_n17309_ & ~new_n17310_;
  assign new_n17312_ = ~new_n4985_ & ~new_n17113_;
  assign new_n17313_ = new_n17113_ & ~new_n17311_;
  assign new_n17314_ = ~new_n17312_ & ~new_n17313_;
  assign new_n17315_ = new_n5051_ & ~new_n17308_;
  assign new_n17316_ = new_n17308_ & ~new_n17314_;
  assign li0674 = new_n17315_ | new_n17316_;
  assign new_n17318_ = lo0789 & new_n17097_;
  assign new_n17319_ = lo0876 & new_n17093_;
  assign new_n17320_ = ~new_n17318_ & ~new_n17319_;
  assign new_n17321_ = lo0803 & new_n17098_;
  assign new_n17322_ = lo0748 & new_n17079_;
  assign new_n17323_ = lo0623 & new_n17080_;
  assign new_n17324_ = ~new_n17322_ & ~new_n17323_;
  assign new_n17325_ = lo0730 & new_n17086_;
  assign new_n17326_ = lo0710 & new_n17087_;
  assign new_n17327_ = ~new_n17325_ & ~new_n17326_;
  assign new_n17328_ = new_n17320_ & ~new_n17321_;
  assign new_n17329_ = new_n17324_ & new_n17328_;
  assign new_n17330_ = new_n17327_ & new_n17329_;
  assign new_n17331_ = lo0296 & ~new_n17105_;
  assign new_n17332_ = lo0199 & lo1031;
  assign new_n17333_ = ~new_n17331_ & ~new_n17332_;
  assign new_n17334_ = ~new_n4765_ & ~new_n17113_;
  assign new_n17335_ = new_n17113_ & ~new_n17333_;
  assign new_n17336_ = ~new_n17334_ & ~new_n17335_;
  assign new_n17337_ = new_n5051_ & ~new_n17330_;
  assign new_n17338_ = new_n17330_ & ~new_n17336_;
  assign li0675 = new_n17337_ | new_n17338_;
  assign new_n17340_ = lo0787 & new_n17097_;
  assign new_n17341_ = lo0881 & new_n17093_;
  assign new_n17342_ = ~new_n17340_ & ~new_n17341_;
  assign new_n17343_ = lo0812 & new_n17098_;
  assign new_n17344_ = lo0746 & new_n17079_;
  assign new_n17345_ = lo0606 & new_n17080_;
  assign new_n17346_ = ~new_n17344_ & ~new_n17345_;
  assign new_n17347_ = lo0729 & new_n17086_;
  assign new_n17348_ = lo0643 & new_n17087_;
  assign new_n17349_ = ~new_n17347_ & ~new_n17348_;
  assign new_n17350_ = new_n17342_ & ~new_n17343_;
  assign new_n17351_ = new_n17346_ & new_n17350_;
  assign new_n17352_ = new_n17349_ & new_n17351_;
  assign new_n17353_ = lo0293 & ~new_n17105_;
  assign new_n17354_ = lo0199 & lo1053;
  assign new_n17355_ = ~new_n17353_ & ~new_n17354_;
  assign new_n17356_ = ~new_n4728_ & ~new_n17113_;
  assign new_n17357_ = new_n17113_ & ~new_n17355_;
  assign new_n17358_ = ~new_n17356_ & ~new_n17357_;
  assign new_n17359_ = new_n5051_ & ~new_n17352_;
  assign new_n17360_ = new_n17352_ & ~new_n17358_;
  assign li0676 = new_n17359_ | new_n17360_;
  assign new_n17362_ = lo0704 & new_n17086_;
  assign new_n17363_ = lo0635 & new_n17087_;
  assign new_n17364_ = ~new_n17362_ & ~new_n17363_;
  assign new_n17365_ = lo0742 & new_n17079_;
  assign new_n17366_ = lo0620 & new_n17080_;
  assign new_n17367_ = lo0870 & new_n17093_;
  assign new_n17368_ = ~new_n17366_ & ~new_n17367_;
  assign new_n17369_ = new_n17364_ & ~new_n17365_;
  assign new_n17370_ = new_n17368_ & new_n17369_;
  assign new_n17371_ = lo0259 & ~new_n17105_;
  assign new_n17372_ = lo0199 & lo1063;
  assign new_n17373_ = ~new_n17371_ & ~new_n17372_;
  assign new_n17374_ = ~new_n5029_ & ~new_n17113_;
  assign new_n17375_ = new_n17113_ & ~new_n17373_;
  assign new_n17376_ = ~new_n17374_ & ~new_n17375_;
  assign new_n17377_ = new_n5051_ & ~new_n17370_;
  assign new_n17378_ = new_n17370_ & ~new_n17376_;
  assign li0677 = new_n17377_ | new_n17378_;
  assign new_n17380_ = lo0688 & new_n17086_;
  assign new_n17381_ = lo0632 & new_n17087_;
  assign new_n17382_ = ~new_n17380_ & ~new_n17381_;
  assign new_n17383_ = lo0760 & new_n17079_;
  assign new_n17384_ = lo0613 & new_n17080_;
  assign new_n17385_ = lo0856 & new_n17093_;
  assign new_n17386_ = ~new_n17384_ & ~new_n17385_;
  assign new_n17387_ = new_n17382_ & ~new_n17383_;
  assign new_n17388_ = new_n17386_ & new_n17387_;
  assign new_n17389_ = lo0260 & ~new_n17105_;
  assign new_n17390_ = lo0199 & lo1061;
  assign new_n17391_ = ~new_n17389_ & ~new_n17390_;
  assign new_n17392_ = ~new_n5005_ & ~new_n17113_;
  assign new_n17393_ = new_n17113_ & ~new_n17391_;
  assign new_n17394_ = ~new_n17392_ & ~new_n17393_;
  assign new_n17395_ = new_n5051_ & ~new_n17388_;
  assign new_n17396_ = new_n17388_ & ~new_n17394_;
  assign li0678 = new_n17395_ | new_n17396_;
  assign new_n17398_ = lo0739 & new_n17079_;
  assign new_n17399_ = lo0621 & new_n17080_;
  assign new_n17400_ = ~new_n17398_ & ~new_n17399_;
  assign new_n17401_ = lo0690 & new_n17086_;
  assign new_n17402_ = lo0665 & new_n17087_;
  assign new_n17403_ = ~new_n17401_ & ~new_n17402_;
  assign new_n17404_ = lo0874 & new_n17093_;
  assign new_n17405_ = lo0791 & new_n17097_;
  assign new_n17406_ = lo0810 & new_n17098_;
  assign new_n17407_ = ~new_n17405_ & ~new_n17406_;
  assign new_n17408_ = new_n17400_ & new_n17403_;
  assign new_n17409_ = ~new_n17404_ & new_n17408_;
  assign new_n17410_ = new_n17407_ & new_n17409_;
  assign new_n17411_ = lo0255 & ~new_n17105_;
  assign new_n17412_ = lo0199 & lo1030;
  assign new_n17413_ = ~new_n17411_ & ~new_n17412_;
  assign new_n17414_ = ~new_n5012_ & ~new_n17113_;
  assign new_n17415_ = new_n17113_ & ~new_n17413_;
  assign new_n17416_ = ~new_n17414_ & ~new_n17415_;
  assign new_n17417_ = new_n5051_ & ~new_n17410_;
  assign new_n17418_ = new_n17410_ & ~new_n17416_;
  assign li0679 = new_n17417_ | new_n17418_;
  assign new_n17420_ = lo0680 & ~li0797;
  assign new_n17421_ = pi011 & li0797;
  assign new_n17422_ = ~new_n17420_ & ~new_n17421_;
  assign li0680 = ~lo0962 & ~new_n17422_;
  assign new_n17424_ = lo0681 & ~li0797;
  assign new_n17425_ = pi014 & li0797;
  assign new_n17426_ = ~new_n17424_ & ~new_n17425_;
  assign li0681 = ~lo0962 & ~new_n17426_;
  assign new_n17428_ = lo0686 & new_n17086_;
  assign new_n17429_ = lo0631 & new_n17087_;
  assign new_n17430_ = ~new_n17428_ & ~new_n17429_;
  assign new_n17431_ = lo0757 & new_n17079_;
  assign new_n17432_ = lo0610 & new_n17080_;
  assign new_n17433_ = lo0848 & new_n17093_;
  assign new_n17434_ = ~new_n17432_ & ~new_n17433_;
  assign new_n17435_ = new_n17430_ & ~new_n17431_;
  assign new_n17436_ = new_n17434_ & new_n17435_;
  assign new_n17437_ = lo0251 & ~new_n17105_;
  assign new_n17438_ = lo0199 & lo1033;
  assign new_n17439_ = ~new_n17437_ & ~new_n17438_;
  assign new_n17440_ = ~new_n4975_ & ~new_n17113_;
  assign new_n17441_ = new_n17113_ & ~new_n17439_;
  assign new_n17442_ = ~new_n17440_ & ~new_n17441_;
  assign new_n17443_ = new_n5051_ & ~new_n17436_;
  assign new_n17444_ = new_n17436_ & ~new_n17442_;
  assign li0682 = new_n17443_ | new_n17444_;
  assign li0823 = lo0953 & new_n16913_;
  assign new_n17447_ = lo0684 & ~li0823;
  assign new_n17448_ = pi041 & li0823;
  assign new_n17449_ = ~new_n17447_ & ~new_n17448_;
  assign li0684 = ~lo0962 & ~new_n17449_;
  assign new_n17451_ = lo0652 & new_n17080_;
  assign new_n17452_ = lo0860 & new_n17093_;
  assign new_n17453_ = ~new_n17451_ & ~new_n17452_;
  assign new_n17454_ = lo0813 & new_n17098_;
  assign new_n17455_ = lo0744 & new_n17079_;
  assign new_n17456_ = lo0728 & new_n17086_;
  assign new_n17457_ = lo0657 & new_n17087_;
  assign new_n17458_ = ~new_n17456_ & ~new_n17457_;
  assign new_n17459_ = new_n17453_ & ~new_n17454_;
  assign new_n17460_ = ~new_n17455_ & new_n17459_;
  assign new_n17461_ = new_n17458_ & new_n17460_;
  assign new_n17462_ = lo1038 & new_n14883_;
  assign new_n17463_ = lo1061 & new_n14878_;
  assign new_n17464_ = lo0199 & lo1070;
  assign new_n17465_ = ~new_n17463_ & ~new_n17464_;
  assign new_n17466_ = ~new_n17462_ & new_n17465_;
  assign new_n17467_ = ~new_n17113_ & ~new_n17466_;
  assign new_n17468_ = ~new_n4917_ & new_n17466_;
  assign new_n17469_ = ~new_n17467_ & ~new_n17468_;
  assign new_n17470_ = new_n5051_ & ~new_n17461_;
  assign new_n17471_ = new_n17461_ & ~new_n17469_;
  assign li0685 = new_n17470_ | new_n17471_;
  assign new_n17473_ = lo0686 & ~li0823;
  assign new_n17474_ = pi024 & li0823;
  assign new_n17475_ = ~new_n17473_ & ~new_n17474_;
  assign li0686 = ~lo0962 & ~new_n17475_;
  assign new_n17477_ = lo0687 & ~li0823;
  assign new_n17478_ = pi038 & li0823;
  assign new_n17479_ = ~new_n17477_ & ~new_n17478_;
  assign li0687 = ~lo0962 & ~new_n17479_;
  assign new_n17481_ = lo0688 & ~li0823;
  assign new_n17482_ = pi026 & li0823;
  assign new_n17483_ = ~new_n17481_ & ~new_n17482_;
  assign li0688 = ~lo0962 & ~new_n17483_;
  assign new_n17485_ = lo0703 & new_n17086_;
  assign new_n17486_ = lo0655 & new_n17087_;
  assign new_n17487_ = ~new_n17485_ & ~new_n17486_;
  assign new_n17488_ = lo0752 & new_n17079_;
  assign new_n17489_ = lo0843 & new_n17093_;
  assign new_n17490_ = lo0658 & new_n17080_;
  assign new_n17491_ = lo0798 & new_n17098_;
  assign new_n17492_ = ~new_n17490_ & ~new_n17491_;
  assign new_n17493_ = new_n17487_ & ~new_n17488_;
  assign new_n17494_ = ~new_n17489_ & new_n17493_;
  assign new_n17495_ = new_n17492_ & new_n17494_;
  assign new_n17496_ = lo1030 & new_n14878_;
  assign new_n17497_ = lo1043 & new_n14883_;
  assign new_n17498_ = lo0199 & lo1073;
  assign new_n17499_ = ~new_n17497_ & ~new_n17498_;
  assign new_n17500_ = ~new_n17496_ & new_n17499_;
  assign new_n17501_ = ~new_n17113_ & ~new_n17500_;
  assign new_n17502_ = ~new_n4924_ & new_n17500_;
  assign new_n17503_ = ~new_n17501_ & ~new_n17502_;
  assign new_n17504_ = new_n5051_ & ~new_n17495_;
  assign new_n17505_ = new_n17495_ & ~new_n17503_;
  assign li0689 = new_n17504_ | new_n17505_;
  assign new_n17507_ = lo0690 & ~li0823;
  assign new_n17508_ = pi019 & li0823;
  assign new_n17509_ = ~new_n17507_ & ~new_n17508_;
  assign li0690 = ~lo0962 & ~new_n17509_;
  assign new_n17511_ = lo0691 & ~li0823;
  assign new_n17512_ = pi018 & li0823;
  assign new_n17513_ = ~new_n17511_ & ~new_n17512_;
  assign li0691 = ~lo0962 & ~new_n17513_;
  assign new_n17515_ = lo0726 & new_n17086_;
  assign new_n17516_ = lo0649 & new_n17087_;
  assign new_n17517_ = ~new_n17515_ & ~new_n17516_;
  assign new_n17518_ = lo0770 & new_n17079_;
  assign new_n17519_ = lo0844 & new_n17093_;
  assign new_n17520_ = lo0656 & new_n17080_;
  assign new_n17521_ = lo0801 & new_n17098_;
  assign new_n17522_ = ~new_n17520_ & ~new_n17521_;
  assign new_n17523_ = new_n17517_ & ~new_n17518_;
  assign new_n17524_ = ~new_n17519_ & new_n17523_;
  assign new_n17525_ = new_n17522_ & new_n17524_;
  assign new_n17526_ = lo1078 & new_n14883_;
  assign new_n17527_ = lo1059 & new_n14878_;
  assign new_n17528_ = lo0199 & lo1072;
  assign new_n17529_ = ~new_n17527_ & ~new_n17528_;
  assign new_n17530_ = ~new_n17526_ & new_n17529_;
  assign new_n17531_ = ~new_n17113_ & ~new_n17530_;
  assign new_n17532_ = ~new_n4934_ & new_n17530_;
  assign new_n17533_ = ~new_n17531_ & ~new_n17532_;
  assign new_n17534_ = new_n5051_ & ~new_n17525_;
  assign new_n17535_ = new_n17525_ & ~new_n17533_;
  assign li0692 = new_n17534_ | new_n17535_;
  assign new_n17537_ = lo0693 & ~li0797;
  assign new_n17538_ = pi040 & li0797;
  assign new_n17539_ = ~new_n17537_ & ~new_n17538_;
  assign li0693 = ~lo0962 & ~new_n17539_;
  assign new_n17541_ = lo0694 & ~li0823;
  assign new_n17542_ = pi039 & li0823;
  assign new_n17543_ = ~new_n17541_ & ~new_n17542_;
  assign li0694 = ~lo0962 & ~new_n17543_;
  assign new_n17545_ = lo0695 & ~li0797;
  assign new_n17546_ = pi022 & li0797;
  assign new_n17547_ = ~new_n17545_ & ~new_n17546_;
  assign li0695 = ~lo0962 & ~new_n17547_;
  assign new_n17549_ = lo0696 & ~li0823;
  assign new_n17550_ = pi011 & li0823;
  assign new_n17551_ = ~new_n17549_ & ~new_n17550_;
  assign li0696 = ~lo0962 & ~new_n17551_;
  assign new_n17553_ = lo0697 & ~li0823;
  assign new_n17554_ = pi040 & li0823;
  assign new_n17555_ = ~new_n17553_ & ~new_n17554_;
  assign li0697 = ~lo0962 & ~new_n17555_;
  assign new_n17557_ = lo0698 & ~li0823;
  assign new_n17558_ = pi027 & li0823;
  assign new_n17559_ = ~new_n17557_ & ~new_n17558_;
  assign li0698 = ~lo0962 & ~new_n17559_;
  assign new_n17561_ = lo0699 & ~li0823;
  assign new_n17562_ = pi014 & li0823;
  assign new_n17563_ = ~new_n17561_ & ~new_n17562_;
  assign li0699 = ~lo0962 & ~new_n17563_;
  assign new_n17565_ = lo0700 & ~li0823;
  assign new_n17566_ = pi021 & li0823;
  assign new_n17567_ = ~new_n17565_ & ~new_n17566_;
  assign li0700 = ~lo0962 & ~new_n17567_;
  assign new_n17569_ = lo0701 & ~li0823;
  assign new_n17570_ = pi034 & li0823;
  assign new_n17571_ = ~new_n17569_ & ~new_n17570_;
  assign li0701 = ~lo0962 & ~new_n17571_;
  assign new_n17573_ = lo0702 & ~li0823;
  assign new_n17574_ = pi028 & li0823;
  assign new_n17575_ = ~new_n17573_ & ~new_n17574_;
  assign li0702 = ~lo0962 & ~new_n17575_;
  assign new_n17577_ = lo0703 & ~li0823;
  assign new_n17578_ = pi035 & li0823;
  assign new_n17579_ = ~new_n17577_ & ~new_n17578_;
  assign li0703 = ~lo0962 & ~new_n17579_;
  assign new_n17581_ = lo0704 & ~li0823;
  assign new_n17582_ = pi023 & li0823;
  assign new_n17583_ = ~new_n17581_ & ~new_n17582_;
  assign li0704 = ~lo0962 & ~new_n17583_;
  assign new_n17585_ = lo0705 & ~li0823;
  assign new_n17586_ = pi036 & li0823;
  assign new_n17587_ = ~new_n17585_ & ~new_n17586_;
  assign li0705 = ~lo0962 & ~new_n17587_;
  assign new_n17589_ = lo0706 & ~li0823;
  assign new_n17590_ = pi016 & li0823;
  assign new_n17591_ = ~new_n17589_ & ~new_n17590_;
  assign li0706 = ~lo0962 & ~new_n17591_;
  assign new_n17593_ = lo0702 & new_n17086_;
  assign new_n17594_ = lo0627 & new_n17087_;
  assign new_n17595_ = ~new_n17593_ & ~new_n17594_;
  assign new_n17596_ = lo0753 & new_n17079_;
  assign new_n17597_ = lo0618 & new_n17080_;
  assign new_n17598_ = lo0847 & new_n17093_;
  assign new_n17599_ = ~new_n17597_ & ~new_n17598_;
  assign new_n17600_ = new_n17595_ & ~new_n17596_;
  assign new_n17601_ = new_n17599_ & new_n17600_;
  assign new_n17602_ = lo1042 & new_n14878_;
  assign new_n17603_ = lo0304 & new_n14883_;
  assign new_n17604_ = lo0199 & lo1049;
  assign new_n17605_ = ~new_n17603_ & ~new_n17604_;
  assign new_n17606_ = ~new_n17602_ & new_n17605_;
  assign new_n17607_ = ~new_n17113_ & ~new_n17606_;
  assign new_n17608_ = ~new_n4809_ & new_n17606_;
  assign new_n17609_ = ~new_n17607_ & ~new_n17608_;
  assign new_n17610_ = new_n5051_ & ~new_n17601_;
  assign new_n17611_ = new_n17601_ & ~new_n17609_;
  assign li0707 = new_n17610_ | new_n17611_;
  assign new_n17613_ = lo0709 & new_n17086_;
  assign new_n17614_ = lo0660 & new_n17087_;
  assign new_n17615_ = ~new_n17613_ & ~new_n17614_;
  assign new_n17616_ = lo0754 & new_n17079_;
  assign new_n17617_ = lo0609 & new_n17080_;
  assign new_n17618_ = lo0857 & new_n17093_;
  assign new_n17619_ = ~new_n17617_ & ~new_n17618_;
  assign new_n17620_ = new_n17615_ & ~new_n17616_;
  assign new_n17621_ = new_n17619_ & new_n17620_;
  assign new_n17622_ = lo1078 & new_n14878_;
  assign new_n17623_ = lo0305 & new_n14883_;
  assign new_n17624_ = lo0199 & lo1052;
  assign new_n17625_ = ~new_n17623_ & ~new_n17624_;
  assign new_n17626_ = ~new_n17622_ & new_n17625_;
  assign new_n17627_ = ~new_n17113_ & ~new_n17626_;
  assign new_n17628_ = ~new_n4846_ & new_n17626_;
  assign new_n17629_ = ~new_n17627_ & ~new_n17628_;
  assign new_n17630_ = new_n5051_ & ~new_n17621_;
  assign new_n17631_ = new_n17621_ & ~new_n17629_;
  assign li0708 = new_n17630_ | new_n17631_;
  assign new_n17633_ = lo0709 & ~li0823;
  assign new_n17634_ = pi029 & li0823;
  assign new_n17635_ = ~new_n17633_ & ~new_n17634_;
  assign li0709 = ~lo0962 & ~new_n17635_;
  assign new_n17637_ = lo0710 & ~li0797;
  assign new_n17638_ = pi017 & li0797;
  assign new_n17639_ = ~new_n17637_ & ~new_n17638_;
  assign li0710 = ~lo0962 & ~new_n17639_;
  assign new_n17641_ = lo0725 & new_n17086_;
  assign new_n17642_ = lo0647 & new_n17087_;
  assign new_n17643_ = ~new_n17641_ & ~new_n17642_;
  assign new_n17644_ = lo0755 & new_n17079_;
  assign new_n17645_ = lo0630 & new_n17080_;
  assign new_n17646_ = lo0858 & new_n17093_;
  assign new_n17647_ = ~new_n17645_ & ~new_n17646_;
  assign new_n17648_ = new_n17643_ & ~new_n17644_;
  assign new_n17649_ = new_n17647_ & new_n17648_;
  assign new_n17650_ = lo1053 & new_n14878_;
  assign new_n17651_ = lo0306 & new_n14883_;
  assign new_n17652_ = lo0199 & lo1081;
  assign new_n17653_ = ~new_n17651_ & ~new_n17652_;
  assign new_n17654_ = ~new_n17650_ & new_n17653_;
  assign new_n17655_ = ~new_n17113_ & ~new_n17654_;
  assign new_n17656_ = ~new_n4853_ & new_n17654_;
  assign new_n17657_ = ~new_n17655_ & ~new_n17656_;
  assign new_n17658_ = new_n5051_ & ~new_n17649_;
  assign new_n17659_ = new_n17649_ & ~new_n17657_;
  assign li0711 = new_n17658_ | new_n17659_;
  assign new_n17661_ = lo0701 & new_n17086_;
  assign new_n17662_ = lo0715 & new_n17087_;
  assign new_n17663_ = ~new_n17661_ & ~new_n17662_;
  assign new_n17664_ = lo0751 & new_n17079_;
  assign new_n17665_ = lo0644 & new_n17080_;
  assign new_n17666_ = lo0842 & new_n17093_;
  assign new_n17667_ = ~new_n17665_ & ~new_n17666_;
  assign new_n17668_ = new_n17663_ & ~new_n17664_;
  assign new_n17669_ = new_n17667_ & new_n17668_;
  assign new_n17670_ = lo1038 & new_n14878_;
  assign new_n17671_ = lo0298 & new_n14883_;
  assign new_n17672_ = lo0199 & lo1029;
  assign new_n17673_ = ~new_n17671_ & ~new_n17672_;
  assign new_n17674_ = ~new_n17670_ & new_n17673_;
  assign new_n17675_ = ~new_n17113_ & ~new_n17674_;
  assign new_n17676_ = ~new_n4829_ & new_n17674_;
  assign new_n17677_ = ~new_n17675_ & ~new_n17676_;
  assign new_n17678_ = new_n5051_ & ~new_n17669_;
  assign new_n17679_ = new_n17669_ & ~new_n17677_;
  assign li0712 = new_n17678_ | new_n17679_;
  assign new_n17681_ = lo0734 & new_n17086_;
  assign new_n17682_ = lo0628 & new_n17087_;
  assign new_n17683_ = ~new_n17681_ & ~new_n17682_;
  assign new_n17684_ = lo0756 & new_n17079_;
  assign new_n17685_ = lo0629 & new_n17080_;
  assign new_n17686_ = lo0854 & new_n17093_;
  assign new_n17687_ = ~new_n17685_ & ~new_n17686_;
  assign new_n17688_ = new_n17683_ & ~new_n17684_;
  assign new_n17689_ = new_n17687_ & new_n17688_;
  assign new_n17690_ = lo1066 & new_n14878_;
  assign new_n17691_ = lo0309 & new_n14883_;
  assign new_n17692_ = lo0199 & lo1045;
  assign new_n17693_ = ~new_n17691_ & ~new_n17692_;
  assign new_n17694_ = ~new_n17690_ & new_n17693_;
  assign new_n17695_ = ~new_n17113_ & ~new_n17694_;
  assign new_n17696_ = ~new_n4792_ & new_n17694_;
  assign new_n17697_ = ~new_n17695_ & ~new_n17696_;
  assign new_n17698_ = new_n5051_ & ~new_n17689_;
  assign new_n17699_ = new_n17689_ & ~new_n17697_;
  assign li0713 = new_n17698_ | new_n17699_;
  assign new_n17701_ = lo0697 & new_n17086_;
  assign new_n17702_ = lo0693 & new_n17087_;
  assign new_n17703_ = ~new_n17701_ & ~new_n17702_;
  assign new_n17704_ = lo0762 & new_n17079_;
  assign new_n17705_ = lo0867 & new_n17093_;
  assign new_n17706_ = lo0653 & new_n17080_;
  assign new_n17707_ = lo0816 & new_n17098_;
  assign new_n17708_ = ~new_n17706_ & ~new_n17707_;
  assign new_n17709_ = new_n17703_ & ~new_n17704_;
  assign new_n17710_ = ~new_n17705_ & new_n17709_;
  assign new_n17711_ = new_n17708_ & new_n17710_;
  assign new_n17712_ = lo1047 & new_n14883_;
  assign new_n17713_ = lo1033 & new_n14878_;
  assign new_n17714_ = lo0199 & lo1051;
  assign new_n17715_ = ~new_n17713_ & ~new_n17714_;
  assign new_n17716_ = ~new_n17712_ & new_n17715_;
  assign new_n17717_ = ~new_n17113_ & ~new_n17716_;
  assign new_n17718_ = ~new_n4897_ & new_n17716_;
  assign new_n17719_ = ~new_n17717_ & ~new_n17718_;
  assign new_n17720_ = new_n5051_ & ~new_n17711_;
  assign new_n17721_ = new_n17711_ & ~new_n17719_;
  assign li0714 = new_n17720_ | new_n17721_;
  assign new_n17723_ = lo0715 & ~li0797;
  assign new_n17724_ = pi034 & li0797;
  assign new_n17725_ = ~new_n17723_ & ~new_n17724_;
  assign li0715 = ~lo0962 & ~new_n17725_;
  assign new_n17727_ = lo0738 & new_n17086_;
  assign new_n17728_ = lo0641 & new_n17087_;
  assign new_n17729_ = ~new_n17727_ & ~new_n17728_;
  assign new_n17730_ = lo0761 & new_n17079_;
  assign new_n17731_ = lo0626 & new_n17080_;
  assign new_n17732_ = lo0845 & new_n17093_;
  assign new_n17733_ = ~new_n17731_ & ~new_n17732_;
  assign new_n17734_ = new_n17729_ & ~new_n17730_;
  assign new_n17735_ = new_n17733_ & new_n17734_;
  assign new_n17736_ = lo1047 & new_n14878_;
  assign new_n17737_ = lo0307 & new_n14883_;
  assign new_n17738_ = lo0199 & lo1037;
  assign new_n17739_ = ~new_n17737_ & ~new_n17738_;
  assign new_n17740_ = ~new_n17736_ & new_n17739_;
  assign new_n17741_ = ~new_n17113_ & ~new_n17740_;
  assign new_n17742_ = ~new_n4799_ & new_n17740_;
  assign new_n17743_ = ~new_n17741_ & ~new_n17742_;
  assign new_n17744_ = new_n5051_ & ~new_n17735_;
  assign new_n17745_ = new_n17735_ & ~new_n17743_;
  assign li0716 = new_n17744_ | new_n17745_;
  assign new_n17747_ = lo0705 & new_n17086_;
  assign new_n17748_ = lo0669 & new_n17087_;
  assign new_n17749_ = ~new_n17747_ & ~new_n17748_;
  assign new_n17750_ = lo0768 & new_n17079_;
  assign new_n17751_ = lo0839 & new_n17093_;
  assign new_n17752_ = lo0645 & new_n17080_;
  assign new_n17753_ = lo0800 & new_n17098_;
  assign new_n17754_ = ~new_n17752_ & ~new_n17753_;
  assign new_n17755_ = new_n17749_ & ~new_n17750_;
  assign new_n17756_ = ~new_n17751_ & new_n17755_;
  assign new_n17757_ = new_n17754_ & new_n17756_;
  assign new_n17758_ = lo1064 & new_n14878_;
  assign new_n17759_ = lo1042 & new_n14883_;
  assign new_n17760_ = lo0199 & lo1068;
  assign new_n17761_ = ~new_n17759_ & ~new_n17760_;
  assign new_n17762_ = ~new_n17758_ & new_n17761_;
  assign new_n17763_ = ~new_n17113_ & ~new_n17762_;
  assign new_n17764_ = ~new_n4880_ & new_n17762_;
  assign new_n17765_ = ~new_n17763_ & ~new_n17764_;
  assign new_n17766_ = new_n5051_ & ~new_n17757_;
  assign new_n17767_ = new_n17757_ & ~new_n17765_;
  assign li0717 = new_n17766_ | new_n17767_;
  assign new_n17769_ = lo0698 & new_n17086_;
  assign new_n17770_ = lo0625 & new_n17087_;
  assign new_n17771_ = ~new_n17769_ & ~new_n17770_;
  assign new_n17772_ = lo0767 & new_n17079_;
  assign new_n17773_ = lo0608 & new_n17080_;
  assign new_n17774_ = lo0853 & new_n17093_;
  assign new_n17775_ = ~new_n17773_ & ~new_n17774_;
  assign new_n17776_ = new_n17771_ & ~new_n17772_;
  assign new_n17777_ = new_n17775_ & new_n17776_;
  assign new_n17778_ = lo1043 & new_n14878_;
  assign new_n17779_ = lo0303 & new_n14883_;
  assign new_n17780_ = lo0199 & lo1074;
  assign new_n17781_ = ~new_n17779_ & ~new_n17780_;
  assign new_n17782_ = ~new_n17778_ & new_n17781_;
  assign new_n17783_ = ~new_n17113_ & ~new_n17782_;
  assign new_n17784_ = ~new_n4836_ & new_n17782_;
  assign new_n17785_ = ~new_n17783_ & ~new_n17784_;
  assign new_n17786_ = new_n5051_ & ~new_n17777_;
  assign new_n17787_ = new_n17777_ & ~new_n17785_;
  assign li0718 = new_n17786_ | new_n17787_;
  assign new_n17789_ = lo0687 & new_n17086_;
  assign new_n17790_ = lo0650 & new_n17087_;
  assign new_n17791_ = ~new_n17789_ & ~new_n17790_;
  assign new_n17792_ = lo0774 & new_n17079_;
  assign new_n17793_ = lo0868 & new_n17093_;
  assign new_n17794_ = lo0636 & new_n17080_;
  assign new_n17795_ = lo0807 & new_n17098_;
  assign new_n17796_ = ~new_n17794_ & ~new_n17795_;
  assign new_n17797_ = new_n17791_ & ~new_n17792_;
  assign new_n17798_ = ~new_n17793_ & new_n17797_;
  assign new_n17799_ = new_n17796_ & new_n17798_;
  assign new_n17800_ = lo1066 & new_n14883_;
  assign new_n17801_ = lo1056 & new_n14878_;
  assign new_n17802_ = lo0199 & lo1057;
  assign new_n17803_ = ~new_n17801_ & ~new_n17802_;
  assign new_n17804_ = ~new_n17800_ & new_n17803_;
  assign new_n17805_ = ~new_n17113_ & ~new_n17804_;
  assign new_n17806_ = ~new_n4904_ & new_n17804_;
  assign new_n17807_ = ~new_n17805_ & ~new_n17806_;
  assign new_n17808_ = new_n5051_ & ~new_n17799_;
  assign new_n17809_ = new_n17799_ & ~new_n17807_;
  assign li0719 = new_n17808_ | new_n17809_;
  assign new_n17811_ = lo0684 & new_n17086_;
  assign new_n17812_ = lo0654 & new_n17087_;
  assign new_n17813_ = ~new_n17811_ & ~new_n17812_;
  assign new_n17814_ = lo0750 & new_n17079_;
  assign new_n17815_ = lo0880 & new_n17093_;
  assign new_n17816_ = lo0651 & new_n17080_;
  assign new_n17817_ = lo0794 & new_n17098_;
  assign new_n17818_ = ~new_n17816_ & ~new_n17817_;
  assign new_n17819_ = new_n17813_ & ~new_n17814_;
  assign new_n17820_ = ~new_n17815_ & new_n17819_;
  assign new_n17821_ = new_n17818_ & new_n17820_;
  assign new_n17822_ = lo1031 & new_n14883_;
  assign new_n17823_ = lo1034 & new_n14878_;
  assign new_n17824_ = lo0199 & lo1075;
  assign new_n17825_ = ~new_n17823_ & ~new_n17824_;
  assign new_n17826_ = ~new_n17822_ & new_n17825_;
  assign new_n17827_ = ~new_n17113_ & ~new_n17826_;
  assign new_n17828_ = ~new_n4887_ & new_n17826_;
  assign new_n17829_ = ~new_n17827_ & ~new_n17828_;
  assign new_n17830_ = new_n5051_ & ~new_n17821_;
  assign new_n17831_ = new_n17821_ & ~new_n17829_;
  assign li0720 = new_n17830_ | new_n17831_;
  assign new_n17833_ = lo0765 & lo0771;
  assign new_n17834_ = lo0773 & new_n17833_;
  assign new_n17835_ = lo0731 & lo0775;
  assign new_n17836_ = new_n17834_ & new_n17835_;
  assign new_n17837_ = lo0769 & new_n17836_;
  assign new_n17838_ = lo0747 & new_n17837_;
  assign new_n17839_ = ~lo0721 & ~new_n17838_;
  assign new_n17840_ = lo0721 & new_n17838_;
  assign new_n17841_ = ~new_n17839_ & ~new_n17840_;
  assign new_n17842_ = lo0945 & new_n17841_;
  assign new_n17843_ = lo0721 & ~lo0945;
  assign new_n17844_ = ~new_n17842_ & ~new_n17843_;
  assign new_n17845_ = ~lo0795 & ~lo0816;
  assign new_n17846_ = ~lo0794 & ~lo0813;
  assign new_n17847_ = new_n17845_ & new_n17846_;
  assign new_n17848_ = ~lo0798 & ~lo0800;
  assign new_n17849_ = ~lo0801 & ~lo0807;
  assign new_n17850_ = new_n17848_ & new_n17849_;
  assign new_n17851_ = lo0775 & ~lo0816;
  assign new_n17852_ = ~lo0775 & lo0816;
  assign new_n17853_ = ~new_n17851_ & ~new_n17852_;
  assign new_n17854_ = lo0731 & ~lo0795;
  assign new_n17855_ = ~lo0731 & lo0795;
  assign new_n17856_ = ~new_n17854_ & ~new_n17855_;
  assign new_n17857_ = lo0769 & ~lo0794;
  assign new_n17858_ = ~lo0769 & lo0794;
  assign new_n17859_ = ~new_n17857_ & ~new_n17858_;
  assign new_n17860_ = lo0721 & lo0813;
  assign new_n17861_ = ~lo0721 & ~lo0813;
  assign new_n17862_ = ~new_n17860_ & ~new_n17861_;
  assign new_n17863_ = lo0747 & ~lo0807;
  assign new_n17864_ = ~lo0747 & lo0807;
  assign new_n17865_ = ~new_n17863_ & ~new_n17864_;
  assign new_n17866_ = ~lo0765 & lo0798;
  assign new_n17867_ = lo0765 & ~lo0798;
  assign new_n17868_ = ~new_n17866_ & ~new_n17867_;
  assign new_n17869_ = new_n17865_ & new_n17868_;
  assign new_n17870_ = lo0773 & ~lo0801;
  assign new_n17871_ = ~lo0773 & lo0801;
  assign new_n17872_ = ~new_n17870_ & ~new_n17871_;
  assign new_n17873_ = lo0771 & ~lo0800;
  assign new_n17874_ = ~lo0771 & lo0800;
  assign new_n17875_ = ~new_n17873_ & ~new_n17874_;
  assign new_n17876_ = new_n17872_ & new_n17875_;
  assign new_n17877_ = ~new_n17862_ & new_n17869_;
  assign new_n17878_ = new_n17876_ & new_n17877_;
  assign new_n17879_ = new_n17853_ & new_n17856_;
  assign new_n17880_ = new_n17859_ & new_n17879_;
  assign li0821 = new_n17878_ & new_n17880_;
  assign new_n17882_ = new_n17847_ & new_n17850_;
  assign li0806 = li0821 & ~new_n17882_;
  assign li0721 = ~new_n17844_ & ~li0806;
  assign new_n17885_ = lo0694 & new_n17086_;
  assign new_n17886_ = lo0732 & new_n17087_;
  assign new_n17887_ = ~new_n17885_ & ~new_n17886_;
  assign new_n17888_ = lo0776 & new_n17079_;
  assign new_n17889_ = lo0851 & new_n17093_;
  assign new_n17890_ = lo0640 & new_n17080_;
  assign new_n17891_ = lo0795 & new_n17098_;
  assign new_n17892_ = ~new_n17890_ & ~new_n17891_;
  assign new_n17893_ = new_n17887_ & ~new_n17888_;
  assign new_n17894_ = ~new_n17889_ & new_n17893_;
  assign new_n17895_ = new_n17892_ & new_n17894_;
  assign new_n17896_ = lo1053 & new_n14883_;
  assign new_n17897_ = lo1063 & new_n14878_;
  assign new_n17898_ = lo0199 & lo1039;
  assign new_n17899_ = ~new_n17897_ & ~new_n17898_;
  assign new_n17900_ = ~new_n17896_ & new_n17899_;
  assign new_n17901_ = ~new_n17113_ & ~new_n17900_;
  assign new_n17902_ = ~new_n4941_ & new_n17900_;
  assign new_n17903_ = ~new_n17901_ & ~new_n17902_;
  assign new_n17904_ = new_n5051_ & ~new_n17895_;
  assign new_n17905_ = new_n17895_ & ~new_n17903_;
  assign li0722 = new_n17904_ | new_n17905_;
  assign new_n17907_ = lo0723 & ~li0823;
  assign new_n17908_ = pi022 & li0823;
  assign new_n17909_ = ~new_n17907_ & ~new_n17908_;
  assign li0723 = ~lo0962 & ~new_n17909_;
  assign new_n17911_ = lo0724 & ~li0823;
  assign new_n17912_ = pi025 & li0823;
  assign new_n17913_ = ~new_n17911_ & ~new_n17912_;
  assign li0724 = ~lo0962 & ~new_n17913_;
  assign new_n17915_ = lo0725 & ~li0823;
  assign new_n17916_ = pi031 & li0823;
  assign new_n17917_ = ~new_n17915_ & ~new_n17916_;
  assign li0725 = ~lo0962 & ~new_n17917_;
  assign new_n17919_ = lo0726 & ~li0823;
  assign new_n17920_ = pi037 & li0823;
  assign new_n17921_ = ~new_n17919_ & ~new_n17920_;
  assign li0726 = ~lo0962 & ~new_n17921_;
  assign new_n17923_ = lo0727 & ~li0823;
  assign new_n17924_ = pi013 & li0823;
  assign new_n17925_ = ~new_n17923_ & ~new_n17924_;
  assign li0727 = ~lo0962 & ~new_n17925_;
  assign new_n17927_ = lo0728 & ~li0823;
  assign new_n17928_ = pi042 & li0823;
  assign new_n17929_ = ~new_n17927_ & ~new_n17928_;
  assign li0728 = ~lo0962 & ~new_n17929_;
  assign new_n17931_ = lo0729 & ~li0823;
  assign new_n17932_ = pi015 & li0823;
  assign new_n17933_ = ~new_n17931_ & ~new_n17932_;
  assign li0729 = ~lo0962 & ~new_n17933_;
  assign new_n17935_ = lo0730 & ~li0823;
  assign new_n17936_ = pi017 & li0823;
  assign new_n17937_ = ~new_n17935_ & ~new_n17936_;
  assign li0730 = ~lo0962 & ~new_n17937_;
  assign new_n17939_ = lo0747 & new_n17834_;
  assign new_n17940_ = ~lo0731 & ~new_n17939_;
  assign new_n17941_ = lo0731 & new_n17939_;
  assign new_n17942_ = ~new_n17940_ & ~new_n17941_;
  assign new_n17943_ = lo0945 & new_n17942_;
  assign new_n17944_ = lo0731 & ~lo0945;
  assign new_n17945_ = ~new_n17943_ & ~new_n17944_;
  assign li0731 = ~li0806 & ~new_n17945_;
  assign new_n17947_ = lo0732 & ~li0797;
  assign new_n17948_ = pi039 & li0797;
  assign new_n17949_ = ~new_n17947_ & ~new_n17948_;
  assign li0732 = ~lo0962 & ~new_n17949_;
  assign new_n17951_ = lo0737 & new_n17086_;
  assign new_n17952_ = lo0648 & new_n17087_;
  assign new_n17953_ = ~new_n17951_ & ~new_n17952_;
  assign new_n17954_ = lo0777 & new_n17079_;
  assign new_n17955_ = lo0619 & new_n17080_;
  assign new_n17956_ = lo0838 & new_n17093_;
  assign new_n17957_ = ~new_n17955_ & ~new_n17956_;
  assign new_n17958_ = new_n17953_ & ~new_n17954_;
  assign new_n17959_ = new_n17957_ & new_n17958_;
  assign new_n17960_ = lo1031 & new_n14878_;
  assign new_n17961_ = lo0308 & new_n14883_;
  assign new_n17962_ = lo0199 & lo1041;
  assign new_n17963_ = ~new_n17961_ & ~new_n17962_;
  assign new_n17964_ = ~new_n17960_ & new_n17963_;
  assign new_n17965_ = ~new_n17113_ & ~new_n17964_;
  assign new_n17966_ = ~new_n4816_ & new_n17964_;
  assign new_n17967_ = ~new_n17965_ & ~new_n17966_;
  assign new_n17968_ = new_n5051_ & ~new_n17959_;
  assign new_n17969_ = new_n17959_ & ~new_n17967_;
  assign li0733 = new_n17968_ | new_n17969_;
  assign new_n17971_ = lo0734 & ~li0823;
  assign new_n17972_ = pi030 & li0823;
  assign new_n17973_ = ~new_n17971_ & ~new_n17972_;
  assign li0734 = ~lo0962 & ~new_n17973_;
  assign new_n17975_ = lo0735 & ~li0823;
  assign new_n17976_ = pi020 & li0823;
  assign new_n17977_ = ~new_n17975_ & ~new_n17976_;
  assign li0735 = ~lo0962 & ~new_n17977_;
  assign new_n17979_ = lo0736 & ~li0823;
  assign new_n17980_ = pi012 & li0823;
  assign new_n17981_ = ~new_n17979_ & ~new_n17980_;
  assign li0736 = ~lo0962 & ~new_n17981_;
  assign new_n17983_ = lo0737 & ~li0823;
  assign new_n17984_ = pi033 & li0823;
  assign new_n17985_ = ~new_n17983_ & ~new_n17984_;
  assign li0737 = ~lo0962 & ~new_n17985_;
  assign new_n17987_ = lo0738 & ~li0823;
  assign new_n17988_ = pi032 & li0823;
  assign new_n17989_ = ~new_n17987_ & ~new_n17988_;
  assign li0738 = ~lo0962 & ~new_n17989_;
  assign li0831 = lo0952 & new_n16803_;
  assign new_n17992_ = lo0739 & li0831;
  assign new_n17993_ = pi019 & ~lo0739;
  assign new_n17994_ = ~new_n17992_ & ~new_n17993_;
  assign li0739 = lo0966 | ~new_n17994_;
  assign new_n17996_ = lo0741 & li0831;
  assign new_n17997_ = pi025 & ~lo0741;
  assign new_n17998_ = ~new_n17996_ & ~new_n17997_;
  assign li0741 = lo0966 | ~new_n17998_;
  assign new_n18000_ = lo0742 & li0831;
  assign new_n18001_ = pi023 & ~lo0742;
  assign new_n18002_ = ~new_n18000_ & ~new_n18001_;
  assign li0742 = lo0966 | ~new_n18002_;
  assign new_n18004_ = lo0743 & li0831;
  assign new_n18005_ = pi020 & ~lo0743;
  assign new_n18006_ = ~new_n18004_ & ~new_n18005_;
  assign li0743 = lo0966 | ~new_n18006_;
  assign new_n18008_ = lo0744 & li0831;
  assign new_n18009_ = pi042 & ~lo0744;
  assign new_n18010_ = ~new_n18008_ & ~new_n18009_;
  assign li0744 = lo0966 | ~new_n18010_;
  assign new_n18012_ = lo0745 & li0831;
  assign new_n18013_ = pi022 & ~lo0745;
  assign new_n18014_ = ~new_n18012_ & ~new_n18013_;
  assign li0745 = lo0966 | ~new_n18014_;
  assign new_n18016_ = lo0746 & li0831;
  assign new_n18017_ = pi015 & ~lo0746;
  assign new_n18018_ = ~new_n18016_ & ~new_n18017_;
  assign li0746 = lo0966 | ~new_n18018_;
  assign new_n18020_ = ~lo0747 & ~new_n17834_;
  assign new_n18021_ = ~new_n17939_ & ~new_n18020_;
  assign new_n18022_ = lo0945 & new_n18021_;
  assign new_n18023_ = lo0747 & ~lo0945;
  assign new_n18024_ = ~new_n18022_ & ~new_n18023_;
  assign li0747 = ~li0806 & ~new_n18024_;
  assign new_n18026_ = lo0748 & li0831;
  assign new_n18027_ = pi017 & ~lo0748;
  assign new_n18028_ = ~new_n18026_ & ~new_n18027_;
  assign li0748 = lo0966 | ~new_n18028_;
  assign new_n18030_ = lo0749 & li0831;
  assign new_n18031_ = pi016 & ~lo0749;
  assign new_n18032_ = ~new_n18030_ & ~new_n18031_;
  assign li0749 = lo0966 | ~new_n18032_;
  assign new_n18034_ = lo0750 & li0831;
  assign new_n18035_ = pi041 & ~lo0750;
  assign new_n18036_ = ~new_n18034_ & ~new_n18035_;
  assign li0750 = lo0966 | ~new_n18036_;
  assign new_n18038_ = lo0751 & li0831;
  assign new_n18039_ = pi034 & ~lo0751;
  assign new_n18040_ = ~new_n18038_ & ~new_n18039_;
  assign li0751 = lo0966 | ~new_n18040_;
  assign new_n18042_ = lo0752 & li0831;
  assign new_n18043_ = pi035 & ~lo0752;
  assign new_n18044_ = ~new_n18042_ & ~new_n18043_;
  assign li0752 = lo0966 | ~new_n18044_;
  assign new_n18046_ = lo0753 & li0831;
  assign new_n18047_ = pi028 & ~lo0753;
  assign new_n18048_ = ~new_n18046_ & ~new_n18047_;
  assign li0753 = lo0966 | ~new_n18048_;
  assign new_n18050_ = lo0754 & li0831;
  assign new_n18051_ = pi029 & ~lo0754;
  assign new_n18052_ = ~new_n18050_ & ~new_n18051_;
  assign li0754 = lo0966 | ~new_n18052_;
  assign new_n18054_ = lo0755 & li0831;
  assign new_n18055_ = pi031 & ~lo0755;
  assign new_n18056_ = ~new_n18054_ & ~new_n18055_;
  assign li0755 = lo0966 | ~new_n18056_;
  assign new_n18058_ = lo0756 & li0831;
  assign new_n18059_ = pi030 & ~lo0756;
  assign new_n18060_ = ~new_n18058_ & ~new_n18059_;
  assign li0756 = lo0966 | ~new_n18060_;
  assign new_n18062_ = lo0757 & li0831;
  assign new_n18063_ = pi024 & ~lo0757;
  assign new_n18064_ = ~new_n18062_ & ~new_n18063_;
  assign li0757 = lo0966 | ~new_n18064_;
  assign new_n18066_ = lo0758 & li0831;
  assign new_n18067_ = pi012 & ~lo0758;
  assign new_n18068_ = ~new_n18066_ & ~new_n18067_;
  assign li0758 = lo0966 | ~new_n18068_;
  assign new_n18070_ = lo0759 & li0831;
  assign new_n18071_ = pi011 & ~lo0759;
  assign new_n18072_ = ~new_n18070_ & ~new_n18071_;
  assign li0759 = lo0966 | ~new_n18072_;
  assign new_n18074_ = lo0760 & li0831;
  assign new_n18075_ = pi026 & ~lo0760;
  assign new_n18076_ = ~new_n18074_ & ~new_n18075_;
  assign li0760 = lo0966 | ~new_n18076_;
  assign new_n18078_ = lo0761 & li0831;
  assign new_n18079_ = pi032 & ~lo0761;
  assign new_n18080_ = ~new_n18078_ & ~new_n18079_;
  assign li0761 = lo0966 | ~new_n18080_;
  assign new_n18082_ = lo0762 & li0831;
  assign new_n18083_ = pi040 & ~lo0762;
  assign new_n18084_ = ~new_n18082_ & ~new_n18083_;
  assign li0762 = lo0966 | ~new_n18084_;
  assign new_n18086_ = lo0763 & li0831;
  assign new_n18087_ = pi014 & ~lo0763;
  assign new_n18088_ = ~new_n18086_ & ~new_n18087_;
  assign li0763 = lo0966 | ~new_n18088_;
  assign new_n18090_ = lo0764 & li0831;
  assign new_n18091_ = pi018 & ~lo0764;
  assign new_n18092_ = ~new_n18090_ & ~new_n18091_;
  assign li0764 = lo0966 | ~new_n18092_;
  assign new_n18094_ = ~lo0765 & ~lo0945;
  assign new_n18095_ = lo0765 & lo0945;
  assign new_n18096_ = ~new_n18094_ & ~new_n18095_;
  assign li0765 = ~li0806 & new_n18096_;
  assign new_n18098_ = lo0766 & li0831;
  assign new_n18099_ = pi021 & ~lo0766;
  assign new_n18100_ = ~new_n18098_ & ~new_n18099_;
  assign li0766 = lo0966 | ~new_n18100_;
  assign new_n18102_ = lo0767 & li0831;
  assign new_n18103_ = pi027 & ~lo0767;
  assign new_n18104_ = ~new_n18102_ & ~new_n18103_;
  assign li0767 = lo0966 | ~new_n18104_;
  assign new_n18106_ = lo0768 & li0831;
  assign new_n18107_ = pi036 & ~lo0768;
  assign new_n18108_ = ~new_n18106_ & ~new_n18107_;
  assign li0768 = lo0966 | ~new_n18108_;
  assign new_n18110_ = lo0747 & lo0773;
  assign new_n18111_ = new_n17833_ & new_n18110_;
  assign new_n18112_ = new_n17835_ & new_n18111_;
  assign new_n18113_ = ~lo0769 & ~new_n18112_;
  assign new_n18114_ = lo0769 & new_n18112_;
  assign new_n18115_ = ~new_n18113_ & ~new_n18114_;
  assign new_n18116_ = lo0945 & new_n18115_;
  assign new_n18117_ = lo0769 & ~lo0945;
  assign new_n18118_ = ~new_n18116_ & ~new_n18117_;
  assign li0769 = ~li0806 & ~new_n18118_;
  assign new_n18120_ = lo0770 & li0831;
  assign new_n18121_ = pi037 & ~lo0770;
  assign new_n18122_ = ~new_n18120_ & ~new_n18121_;
  assign li0770 = lo0966 | ~new_n18122_;
  assign new_n18124_ = lo0771 & ~lo0945;
  assign new_n18125_ = lo0765 & ~lo0771;
  assign new_n18126_ = ~lo0765 & lo0771;
  assign new_n18127_ = ~new_n18125_ & ~new_n18126_;
  assign new_n18128_ = lo0945 & ~new_n18127_;
  assign new_n18129_ = ~new_n18124_ & ~new_n18128_;
  assign li0771 = ~li0806 & ~new_n18129_;
  assign new_n18131_ = lo0772 & li0831;
  assign new_n18132_ = pi013 & ~lo0772;
  assign new_n18133_ = ~new_n18131_ & ~new_n18132_;
  assign li0772 = lo0966 | ~new_n18133_;
  assign new_n18135_ = ~lo0773 & ~new_n17833_;
  assign new_n18136_ = ~new_n17834_ & ~new_n18135_;
  assign new_n18137_ = lo0945 & new_n18136_;
  assign new_n18138_ = lo0773 & ~lo0945;
  assign new_n18139_ = ~new_n18137_ & ~new_n18138_;
  assign li0773 = ~li0806 & ~new_n18139_;
  assign new_n18141_ = lo0774 & li0831;
  assign new_n18142_ = pi038 & ~lo0774;
  assign new_n18143_ = ~new_n18141_ & ~new_n18142_;
  assign li0774 = lo0966 | ~new_n18143_;
  assign new_n18145_ = lo0771 & new_n18110_;
  assign new_n18146_ = lo0731 & new_n18145_;
  assign new_n18147_ = lo0765 & new_n18146_;
  assign new_n18148_ = ~lo0775 & ~new_n18147_;
  assign new_n18149_ = lo0775 & new_n18147_;
  assign new_n18150_ = ~new_n18148_ & ~new_n18149_;
  assign new_n18151_ = lo0945 & new_n18150_;
  assign new_n18152_ = lo0775 & ~lo0945;
  assign new_n18153_ = ~new_n18151_ & ~new_n18152_;
  assign li0775 = ~li0806 & ~new_n18153_;
  assign new_n18155_ = lo0776 & li0831;
  assign new_n18156_ = pi039 & ~lo0776;
  assign new_n18157_ = ~new_n18155_ & ~new_n18156_;
  assign li0776 = lo0966 | ~new_n18157_;
  assign new_n18159_ = lo0777 & li0831;
  assign new_n18160_ = pi033 & ~lo0777;
  assign new_n18161_ = ~new_n18159_ & ~new_n18160_;
  assign li0777 = lo0966 | ~new_n18161_;
  assign new_n18163_ = ~lo0956 & ~lo1079;
  assign new_n18164_ = lo0832 & new_n18163_;
  assign new_n18165_ = ~lo1040 & ~lo1077;
  assign new_n18166_ = new_n18164_ & new_n18165_;
  assign new_n18167_ = lo0968 & new_n18166_;
  assign new_n18168_ = pi011 & ~new_n18167_;
  assign new_n18169_ = ~pi011 & lo0778;
  assign li0778 = new_n18168_ | new_n18169_;
  assign li0779 = lo0779 | new_n16863_;
  assign li0780 = lo0780 | new_n16768_;
  assign new_n18173_ = pi012 & ~new_n18167_;
  assign new_n18174_ = ~pi012 & lo0781;
  assign li0781 = new_n18173_ | new_n18174_;
  assign new_n18176_ = ~lo0979 & ~lo0984;
  assign new_n18177_ = ~new_n16815_ & ~new_n18176_;
  assign li0782 = new_n16767_ | ~new_n18177_;
  assign new_n18179_ = pi020 & ~new_n18167_;
  assign new_n18180_ = ~pi020 & lo0783;
  assign li0783 = new_n18179_ | new_n18180_;
  assign new_n18182_ = pi021 & ~new_n18167_;
  assign new_n18183_ = ~pi021 & lo0784;
  assign li0784 = new_n18182_ | new_n18183_;
  assign new_n18185_ = pi013 & ~new_n18167_;
  assign new_n18186_ = ~pi013 & lo0785;
  assign li0785 = new_n18185_ | new_n18186_;
  assign new_n18188_ = lo0786 & lo0954;
  assign new_n18189_ = lo0024 & ~lo0954;
  assign li0786 = new_n18188_ | new_n18189_;
  assign new_n18191_ = pi015 & ~new_n18167_;
  assign new_n18192_ = ~pi015 & lo0787;
  assign li0787 = new_n18191_ | new_n18192_;
  assign new_n18194_ = pi016 & ~new_n18167_;
  assign new_n18195_ = ~pi016 & lo0788;
  assign li0788 = new_n18194_ | new_n18195_;
  assign new_n18197_ = pi017 & ~new_n18167_;
  assign new_n18198_ = ~pi017 & lo0789;
  assign li0789 = new_n18197_ | new_n18198_;
  assign new_n18200_ = pi018 & ~new_n18167_;
  assign new_n18201_ = ~pi018 & lo0790;
  assign li0790 = new_n18200_ | new_n18201_;
  assign new_n18203_ = pi019 & ~new_n18167_;
  assign new_n18204_ = ~pi019 & lo0791;
  assign li0791 = new_n18203_ | new_n18204_;
  assign new_n18206_ = pi014 & ~new_n18167_;
  assign new_n18207_ = ~pi014 & lo0792;
  assign li0792 = new_n18206_ | new_n18207_;
  assign new_n18209_ = ~lo0968 & new_n18165_;
  assign new_n18210_ = new_n18164_ & new_n18209_;
  assign new_n18211_ = lo0794 & new_n18210_;
  assign new_n18212_ = pi041 & ~lo0794;
  assign li0794 = new_n18211_ | new_n18212_;
  assign new_n18214_ = lo0795 & new_n18210_;
  assign new_n18215_ = pi039 & ~lo0795;
  assign li0795 = new_n18214_ | new_n18215_;
  assign new_n18217_ = lo0278 & lo0281;
  assign new_n18218_ = lo0266 & lo0279;
  assign new_n18219_ = lo0269 & new_n18218_;
  assign new_n18220_ = lo0280 & new_n18219_;
  assign new_n18221_ = new_n18217_ & new_n18220_;
  assign new_n18222_ = lo0282 & new_n18221_;
  assign new_n18223_ = lo0277 & new_n18222_;
  assign new_n18224_ = lo0270 & new_n18223_;
  assign new_n18225_ = lo0264 & ~new_n18224_;
  assign new_n18226_ = ~lo0264 & new_n18224_;
  assign li0796 = new_n18225_ | new_n18226_;
  assign new_n18228_ = lo0798 & new_n18210_;
  assign new_n18229_ = pi035 & ~lo0798;
  assign li0798 = new_n18228_ | new_n18229_;
  assign new_n18231_ = lo0799 & new_n18210_;
  assign new_n18232_ = pi018 & ~lo0799;
  assign li0799 = new_n18231_ | new_n18232_;
  assign new_n18234_ = lo0800 & new_n18210_;
  assign new_n18235_ = pi036 & ~lo0800;
  assign li0800 = new_n18234_ | new_n18235_;
  assign new_n18237_ = lo0801 & new_n18210_;
  assign new_n18238_ = pi037 & ~lo0801;
  assign li0801 = new_n18237_ | new_n18238_;
  assign new_n18240_ = new_n17053_ & new_n17057_;
  assign new_n18241_ = lo0269 & lo0281;
  assign new_n18242_ = lo0270 & lo0282;
  assign new_n18243_ = new_n18241_ & new_n18242_;
  assign new_n18244_ = new_n18240_ & new_n18243_;
  assign new_n18245_ = lo0274 & new_n18244_;
  assign li0802 = lo0265 & new_n18245_;
  assign new_n18247_ = lo0803 & new_n18210_;
  assign new_n18248_ = pi017 & ~lo0803;
  assign li0803 = new_n18247_ | new_n18248_;
  assign new_n18250_ = lo0804 & new_n18210_;
  assign new_n18251_ = pi020 & ~lo0804;
  assign li0804 = new_n18250_ | new_n18251_;
  assign new_n18253_ = lo0270 & ~new_n17056_;
  assign new_n18254_ = ~lo0270 & new_n17056_;
  assign li0805 = new_n18253_ | new_n18254_;
  assign new_n18256_ = lo0807 & new_n18210_;
  assign new_n18257_ = pi038 & ~lo0807;
  assign li0807 = new_n18256_ | new_n18257_;
  assign new_n18259_ = lo0808 & new_n18210_;
  assign new_n18260_ = pi012 & ~lo0808;
  assign li0808 = new_n18259_ | new_n18260_;
  assign new_n18262_ = lo0809 & new_n18210_;
  assign new_n18263_ = pi014 & ~lo0809;
  assign li0809 = new_n18262_ | new_n18263_;
  assign new_n18265_ = lo0810 & new_n18210_;
  assign new_n18266_ = pi019 & ~lo0810;
  assign li0810 = new_n18265_ | new_n18266_;
  assign new_n18268_ = lo0811 & new_n18210_;
  assign new_n18269_ = pi013 & ~lo0811;
  assign li0811 = new_n18268_ | new_n18269_;
  assign new_n18271_ = lo0812 & new_n18210_;
  assign new_n18272_ = pi015 & ~lo0812;
  assign li0812 = new_n18271_ | new_n18272_;
  assign new_n18274_ = lo0813 & new_n18210_;
  assign new_n18275_ = pi042 & ~lo0813;
  assign li0813 = new_n18274_ | new_n18275_;
  assign new_n18277_ = lo0814 & new_n18210_;
  assign new_n18278_ = pi016 & ~lo0814;
  assign li0814 = new_n18277_ | new_n18278_;
  assign new_n18280_ = lo0815 & new_n18210_;
  assign new_n18281_ = pi021 & ~lo0815;
  assign li0815 = new_n18280_ | new_n18281_;
  assign new_n18283_ = lo0816 & new_n18210_;
  assign new_n18284_ = pi040 & ~lo0816;
  assign li0816 = new_n18283_ | new_n18284_;
  assign new_n18286_ = ~lo0269 & new_n17053_;
  assign new_n18287_ = lo0269 & ~new_n17053_;
  assign li0817 = new_n18286_ | new_n18287_;
  assign new_n18289_ = new_n17057_ & new_n18242_;
  assign new_n18290_ = lo0280 & new_n18241_;
  assign new_n18291_ = new_n17052_ & new_n18290_;
  assign new_n18292_ = new_n18289_ & new_n18291_;
  assign new_n18293_ = ~lo0265 & new_n18292_;
  assign new_n18294_ = lo0265 & ~new_n18292_;
  assign li0819 = new_n18293_ | new_n18294_;
  assign new_n18296_ = new_n17053_ & new_n18243_;
  assign new_n18297_ = ~lo0277 & new_n18296_;
  assign new_n18298_ = lo0277 & ~new_n18296_;
  assign li0820 = new_n18297_ | new_n18298_;
  assign li0822 = ~lo0811 & ~lo0893;
  assign new_n18301_ = new_n3679_ & new_n5051_;
  assign new_n18302_ = pi003 & new_n3677_;
  assign new_n18303_ = ~lo0982 & ~new_n18301_;
  assign li0824 = new_n18302_ & ~new_n18303_;
  assign new_n18305_ = pi038 & ~pi040;
  assign new_n18306_ = ~pi038 & pi040;
  assign new_n18307_ = ~new_n18305_ & ~new_n18306_;
  assign new_n18308_ = pi036 & ~pi041;
  assign new_n18309_ = ~pi036 & pi041;
  assign new_n18310_ = ~new_n18308_ & ~new_n18309_;
  assign new_n18311_ = new_n18307_ & ~new_n18310_;
  assign new_n18312_ = ~new_n18307_ & new_n18310_;
  assign new_n18313_ = ~new_n18311_ & ~new_n18312_;
  assign new_n18314_ = pi037 & ~pi039;
  assign new_n18315_ = ~pi037 & pi039;
  assign new_n18316_ = ~new_n18314_ & ~new_n18315_;
  assign new_n18317_ = pi035 & ~pi042;
  assign new_n18318_ = ~pi035 & pi042;
  assign new_n18319_ = ~new_n18317_ & ~new_n18318_;
  assign new_n18320_ = new_n18316_ & ~new_n18319_;
  assign new_n18321_ = ~new_n18316_ & new_n18319_;
  assign new_n18322_ = ~new_n18320_ & ~new_n18321_;
  assign new_n18323_ = new_n18313_ & ~new_n18322_;
  assign new_n18324_ = ~new_n18313_ & new_n18322_;
  assign new_n18325_ = ~new_n18323_ & ~new_n18324_;
  assign new_n18326_ = ~lo0123 & new_n17112_;
  assign new_n18327_ = ~new_n18325_ & new_n18326_;
  assign new_n18328_ = lo0825 & new_n18325_;
  assign li0825 = new_n18327_ | new_n18328_;
  assign new_n18330_ = pi028 & ~pi033;
  assign new_n18331_ = ~pi028 & pi033;
  assign new_n18332_ = ~new_n18330_ & ~new_n18331_;
  assign new_n18333_ = pi030 & ~pi032;
  assign new_n18334_ = ~pi030 & pi032;
  assign new_n18335_ = ~new_n18333_ & ~new_n18334_;
  assign new_n18336_ = new_n18332_ & ~new_n18335_;
  assign new_n18337_ = ~new_n18332_ & new_n18335_;
  assign new_n18338_ = ~new_n18336_ & ~new_n18337_;
  assign new_n18339_ = pi029 & ~pi031;
  assign new_n18340_ = ~pi029 & pi031;
  assign new_n18341_ = ~new_n18339_ & ~new_n18340_;
  assign new_n18342_ = pi027 & ~pi034;
  assign new_n18343_ = ~pi027 & pi034;
  assign new_n18344_ = ~new_n18342_ & ~new_n18343_;
  assign new_n18345_ = new_n18341_ & ~new_n18344_;
  assign new_n18346_ = ~new_n18341_ & new_n18344_;
  assign new_n18347_ = ~new_n18345_ & ~new_n18346_;
  assign new_n18348_ = new_n18338_ & ~new_n18347_;
  assign new_n18349_ = ~new_n18338_ & new_n18347_;
  assign new_n18350_ = ~new_n18348_ & ~new_n18349_;
  assign new_n18351_ = new_n18326_ & ~new_n18350_;
  assign new_n18352_ = lo0826 & new_n18350_;
  assign li0826 = new_n18351_ | new_n18352_;
  assign new_n18354_ = pi012 & ~pi017;
  assign new_n18355_ = ~pi012 & pi017;
  assign new_n18356_ = ~new_n18354_ & ~new_n18355_;
  assign new_n18357_ = pi014 & ~pi016;
  assign new_n18358_ = ~pi014 & pi016;
  assign new_n18359_ = ~new_n18357_ & ~new_n18358_;
  assign new_n18360_ = new_n18356_ & ~new_n18359_;
  assign new_n18361_ = ~new_n18356_ & new_n18359_;
  assign new_n18362_ = ~new_n18360_ & ~new_n18361_;
  assign new_n18363_ = pi011 & ~pi018;
  assign new_n18364_ = ~pi011 & pi018;
  assign new_n18365_ = ~new_n18363_ & ~new_n18364_;
  assign new_n18366_ = pi013 & ~pi015;
  assign new_n18367_ = ~pi013 & pi015;
  assign new_n18368_ = ~new_n18366_ & ~new_n18367_;
  assign new_n18369_ = new_n18365_ & ~new_n18368_;
  assign new_n18370_ = ~new_n18365_ & new_n18368_;
  assign new_n18371_ = ~new_n18369_ & ~new_n18370_;
  assign new_n18372_ = new_n18362_ & ~new_n18371_;
  assign new_n18373_ = ~new_n18362_ & new_n18371_;
  assign new_n18374_ = ~new_n18372_ & ~new_n18373_;
  assign new_n18375_ = new_n18326_ & ~new_n18374_;
  assign new_n18376_ = lo0827 & new_n18374_;
  assign li0827 = new_n18375_ | new_n18376_;
  assign new_n18378_ = pi022 & ~pi024;
  assign new_n18379_ = ~pi022 & pi024;
  assign new_n18380_ = ~new_n18378_ & ~new_n18379_;
  assign new_n18381_ = pi020 & ~pi025;
  assign new_n18382_ = ~pi020 & pi025;
  assign new_n18383_ = ~new_n18381_ & ~new_n18382_;
  assign new_n18384_ = new_n18380_ & ~new_n18383_;
  assign new_n18385_ = ~new_n18380_ & new_n18383_;
  assign new_n18386_ = ~new_n18384_ & ~new_n18385_;
  assign new_n18387_ = pi021 & ~pi023;
  assign new_n18388_ = ~pi021 & pi023;
  assign new_n18389_ = ~new_n18387_ & ~new_n18388_;
  assign new_n18390_ = pi019 & ~pi026;
  assign new_n18391_ = ~pi019 & pi026;
  assign new_n18392_ = ~new_n18390_ & ~new_n18391_;
  assign new_n18393_ = new_n18389_ & ~new_n18392_;
  assign new_n18394_ = ~new_n18389_ & new_n18392_;
  assign new_n18395_ = ~new_n18393_ & ~new_n18394_;
  assign new_n18396_ = new_n18386_ & ~new_n18395_;
  assign new_n18397_ = ~new_n18386_ & new_n18395_;
  assign new_n18398_ = ~new_n18396_ & ~new_n18397_;
  assign new_n18399_ = new_n18326_ & ~new_n18398_;
  assign new_n18400_ = lo0828 & new_n18398_;
  assign li0828 = new_n18399_ | new_n18400_;
  assign new_n18402_ = new_n4666_ & new_n5051_;
  assign new_n18403_ = ~lo0951 & ~new_n18402_;
  assign li0829 = pi003 & ~new_n18403_;
  assign new_n18405_ = lo0278 & new_n18220_;
  assign new_n18406_ = ~lo0281 & new_n18405_;
  assign new_n18407_ = lo0281 & ~new_n18405_;
  assign li0830 = new_n18406_ | new_n18407_;
  assign new_n18409_ = pi002 & new_n3673_;
  assign new_n18410_ = ~lo0832 & new_n18409_;
  assign li0832 = new_n5055_ & new_n18410_;
  assign new_n18412_ = lo0833 & ~new_n3673_;
  assign li0833 = new_n18409_ | new_n18412_;
  assign li0835 = lo0946 & new_n3673_;
  assign new_n18415_ = ~lo0282 & new_n18291_;
  assign new_n18416_ = lo0282 & ~new_n18291_;
  assign li0836 = new_n18415_ | new_n18416_;
  assign new_n18418_ = ~lo0955 & lo1043;
  assign new_n18419_ = lo0837 & ~lo1043;
  assign li0837 = new_n18418_ | new_n18419_;
  assign new_n18421_ = ~lo0955 & lo1041;
  assign new_n18422_ = lo0838 & ~lo1041;
  assign li0838 = new_n18421_ | new_n18422_;
  assign new_n18424_ = ~lo0955 & lo1068;
  assign new_n18425_ = lo0839 & ~lo1068;
  assign li0839 = new_n18424_ | new_n18425_;
  assign new_n18427_ = lo0840 & new_n3673_;
  assign new_n18428_ = pi107 & ~lo0840;
  assign li0840 = new_n18427_ | new_n18428_;
  assign new_n18430_ = ~lo0955 & lo1029;
  assign new_n18431_ = lo0842 & ~lo1029;
  assign li0842 = new_n18430_ | new_n18431_;
  assign new_n18433_ = ~lo0955 & lo1073;
  assign new_n18434_ = lo0843 & ~lo1073;
  assign li0843 = new_n18433_ | new_n18434_;
  assign new_n18436_ = ~lo0955 & lo1072;
  assign new_n18437_ = lo0844 & ~lo1072;
  assign li0844 = new_n18436_ | new_n18437_;
  assign new_n18439_ = ~lo0955 & lo1037;
  assign new_n18440_ = lo0845 & ~lo1037;
  assign li0845 = new_n18439_ | new_n18440_;
  assign new_n18442_ = pi045 & new_n14975_;
  assign new_n18443_ = ~pi045 & lo0846;
  assign li0846 = new_n18442_ | new_n18443_;
  assign new_n18445_ = ~lo0955 & lo1049;
  assign new_n18446_ = lo0847 & ~lo1049;
  assign li0847 = new_n18445_ | new_n18446_;
  assign new_n18448_ = ~lo0955 & lo1033;
  assign new_n18449_ = lo0848 & ~lo1033;
  assign li0848 = new_n18448_ | new_n18449_;
  assign new_n18451_ = lo0849 & new_n3673_;
  assign new_n18452_ = pi109 & ~lo0849;
  assign li0849 = new_n18451_ | new_n18452_;
  assign new_n18454_ = ~lo0955 & lo1042;
  assign new_n18455_ = lo0850 & ~lo1042;
  assign li0850 = new_n18454_ | new_n18455_;
  assign new_n18457_ = ~lo0955 & lo1039;
  assign new_n18458_ = lo0851 & ~lo1039;
  assign li0851 = new_n18457_ | new_n18458_;
  assign new_n18460_ = ~lo0955 & lo1056;
  assign new_n18461_ = lo0852 & ~lo1056;
  assign li0852 = new_n18460_ | new_n18461_;
  assign new_n18463_ = ~lo0955 & lo1074;
  assign new_n18464_ = lo0853 & ~lo1074;
  assign li0853 = new_n18463_ | new_n18464_;
  assign new_n18466_ = ~lo0955 & lo1045;
  assign new_n18467_ = lo0854 & ~lo1045;
  assign li0854 = new_n18466_ | new_n18467_;
  assign new_n18469_ = ~lo0955 & lo1059;
  assign new_n18470_ = lo0855 & ~lo1059;
  assign li0855 = new_n18469_ | new_n18470_;
  assign new_n18472_ = ~lo0955 & lo1061;
  assign new_n18473_ = lo0856 & ~lo1061;
  assign li0856 = new_n18472_ | new_n18473_;
  assign new_n18475_ = ~lo0955 & lo1052;
  assign new_n18476_ = lo0857 & ~lo1052;
  assign li0857 = new_n18475_ | new_n18476_;
  assign new_n18478_ = ~lo0955 & lo1081;
  assign new_n18479_ = lo0858 & ~lo1081;
  assign li0858 = new_n18478_ | new_n18479_;
  assign new_n18481_ = ~lo0955 & lo1064;
  assign new_n18482_ = lo0859 & ~lo1064;
  assign li0859 = new_n18481_ | new_n18482_;
  assign new_n18484_ = ~lo0955 & lo1070;
  assign new_n18485_ = lo0860 & ~lo1070;
  assign li0860 = new_n18484_ | new_n18485_;
  assign new_n18487_ = pi052 & new_n14975_;
  assign new_n18488_ = ~pi052 & lo0861;
  assign li0861 = new_n18487_ | new_n18488_;
  assign new_n18490_ = pi050 & new_n14975_;
  assign new_n18491_ = ~pi050 & lo0862;
  assign li0862 = new_n18490_ | new_n18491_;
  assign new_n18493_ = lo0863 & new_n3673_;
  assign new_n18494_ = pi110 & ~lo0863;
  assign li0863 = new_n18493_ | new_n18494_;
  assign new_n18496_ = lo0864 & new_n3673_;
  assign new_n18497_ = pi108 & ~lo0864;
  assign li0864 = new_n18496_ | new_n18497_;
  assign new_n18499_ = ~lo0955 & lo1034;
  assign new_n18500_ = lo0865 & ~lo1034;
  assign li0865 = new_n18499_ | new_n18500_;
  assign new_n18502_ = ~lo0955 & lo1047;
  assign new_n18503_ = lo0866 & ~lo1047;
  assign li0866 = new_n18502_ | new_n18503_;
  assign new_n18505_ = ~lo0955 & lo1051;
  assign new_n18506_ = lo0867 & ~lo1051;
  assign li0867 = new_n18505_ | new_n18506_;
  assign new_n18508_ = ~lo0955 & lo1057;
  assign new_n18509_ = lo0868 & ~lo1057;
  assign li0868 = new_n18508_ | new_n18509_;
  assign new_n18511_ = pi051 & new_n14975_;
  assign new_n18512_ = ~pi051 & lo0869;
  assign li0869 = new_n18511_ | new_n18512_;
  assign new_n18514_ = ~lo0955 & lo1063;
  assign new_n18515_ = lo0870 & ~lo1063;
  assign li0870 = new_n18514_ | new_n18515_;
  assign new_n18517_ = ~lo0955 & lo1066;
  assign new_n18518_ = lo0871 & ~lo1066;
  assign li0871 = new_n18517_ | new_n18518_;
  assign new_n18520_ = ~lo0955 & lo1078;
  assign new_n18521_ = lo0872 & ~lo1078;
  assign li0872 = new_n18520_ | new_n18521_;
  assign new_n18523_ = ~lo0955 & lo1038;
  assign new_n18524_ = lo0873 & ~lo1038;
  assign li0873 = new_n18523_ | new_n18524_;
  assign new_n18526_ = ~lo0955 & lo1030;
  assign new_n18527_ = lo0874 & ~lo1030;
  assign li0874 = new_n18526_ | new_n18527_;
  assign new_n18529_ = pi047 & new_n14975_;
  assign new_n18530_ = ~pi047 & lo0875;
  assign li0875 = new_n18529_ | new_n18530_;
  assign new_n18532_ = ~lo0955 & lo1031;
  assign new_n18533_ = lo0876 & ~lo1031;
  assign li0876 = new_n18532_ | new_n18533_;
  assign new_n18535_ = pi049 & new_n14975_;
  assign new_n18536_ = ~pi049 & lo0877;
  assign li0877 = new_n18535_ | new_n18536_;
  assign new_n18538_ = pi048 & new_n14975_;
  assign new_n18539_ = ~pi048 & lo0878;
  assign li0878 = new_n18538_ | new_n18539_;
  assign new_n18541_ = pi046 & new_n14975_;
  assign new_n18542_ = ~pi046 & lo0879;
  assign li0879 = new_n18541_ | new_n18542_;
  assign new_n18544_ = ~lo0955 & lo1075;
  assign new_n18545_ = lo0880 & ~lo1075;
  assign li0880 = new_n18544_ | new_n18545_;
  assign new_n18547_ = ~lo0955 & lo1053;
  assign new_n18548_ = lo0881 & ~lo1053;
  assign li0881 = new_n18547_ | new_n18548_;
  assign new_n18550_ = pi018 & new_n18326_;
  assign new_n18551_ = ~pi018 & lo0883;
  assign li0883 = new_n18550_ | new_n18551_;
  assign new_n18553_ = pi035 & new_n18326_;
  assign new_n18554_ = ~pi035 & lo0884;
  assign li0884 = new_n18553_ | new_n18554_;
  assign new_n18556_ = pi036 & new_n18326_;
  assign new_n18557_ = ~pi036 & lo0885;
  assign li0885 = new_n18556_ | new_n18557_;
  assign new_n18559_ = pi020 & new_n18326_;
  assign new_n18560_ = ~pi020 & lo0886;
  assign li0886 = new_n18559_ | new_n18560_;
  assign new_n18562_ = pi011 & new_n18326_;
  assign new_n18563_ = ~pi011 & lo0887;
  assign li0887 = new_n18562_ | new_n18563_;
  assign new_n18565_ = pi031 & new_n18326_;
  assign new_n18566_ = ~pi031 & lo0888;
  assign li0888 = new_n18565_ | new_n18566_;
  assign new_n18568_ = pi014 & new_n18326_;
  assign new_n18569_ = ~pi014 & lo0889;
  assign li0889 = new_n18568_ | new_n18569_;
  assign new_n18571_ = pi037 & new_n18326_;
  assign new_n18572_ = ~pi037 & lo0890;
  assign li0890 = new_n18571_ | new_n18572_;
  assign new_n18574_ = pi027 & new_n18326_;
  assign new_n18575_ = ~pi027 & lo0891;
  assign li0891 = new_n18574_ | new_n18575_;
  assign new_n18577_ = pi012 & new_n18326_;
  assign new_n18578_ = ~pi012 & lo0892;
  assign li0892 = new_n18577_ | new_n18578_;
  assign new_n18580_ = pi030 & new_n18326_;
  assign new_n18581_ = ~pi030 & lo0894;
  assign li0894 = new_n18580_ | new_n18581_;
  assign new_n18583_ = pi024 & new_n18326_;
  assign new_n18584_ = ~pi024 & lo0895;
  assign li0895 = new_n18583_ | new_n18584_;
  assign new_n18586_ = pi029 & new_n18326_;
  assign new_n18587_ = ~pi029 & lo0896;
  assign li0896 = new_n18586_ | new_n18587_;
  assign new_n18589_ = pi040 & new_n18326_;
  assign new_n18590_ = ~pi040 & lo0898;
  assign li0898 = new_n18589_ | new_n18590_;
  assign new_n18592_ = pi026 & new_n18326_;
  assign new_n18593_ = ~pi026 & lo0899;
  assign li0899 = new_n18592_ | new_n18593_;
  assign new_n18595_ = pi021 & new_n18326_;
  assign new_n18596_ = ~pi021 & lo0900;
  assign li0900 = new_n18595_ | new_n18596_;
  assign new_n18598_ = pi022 & new_n18326_;
  assign new_n18599_ = ~pi022 & lo0902;
  assign li0902 = new_n18598_ | new_n18599_;
  assign new_n18601_ = pi032 & new_n18326_;
  assign new_n18602_ = ~pi032 & lo0903;
  assign li0903 = new_n18601_ | new_n18602_;
  assign new_n18604_ = pi038 & new_n18326_;
  assign new_n18605_ = ~pi038 & lo0904;
  assign li0904 = new_n18604_ | new_n18605_;
  assign new_n18607_ = pi042 & new_n18326_;
  assign new_n18608_ = ~pi042 & lo0905;
  assign li0905 = new_n18607_ | new_n18608_;
  assign new_n18610_ = pi039 & new_n18326_;
  assign new_n18611_ = ~pi039 & lo0906;
  assign li0906 = new_n18610_ | new_n18611_;
  assign new_n18613_ = ~lo0604 & ~lo0979;
  assign new_n18614_ = ~lo0615 & lo0979;
  assign new_n18615_ = ~new_n18613_ & ~new_n18614_;
  assign new_n18616_ = lo0624 & lo0979;
  assign new_n18617_ = lo0598 & ~lo0624;
  assign new_n18618_ = ~new_n18616_ & ~new_n18617_;
  assign new_n18619_ = new_n18615_ & new_n18618_;
  assign new_n18620_ = lo0782 & new_n18619_;
  assign new_n18621_ = ~lo0782 & lo0907;
  assign li0907 = new_n18620_ | new_n18621_;
  assign new_n18623_ = pi033 & new_n18326_;
  assign new_n18624_ = ~pi033 & lo0908;
  assign li0908 = new_n18623_ | new_n18624_;
  assign new_n18626_ = pi016 & new_n18326_;
  assign new_n18627_ = ~pi016 & lo0909;
  assign li0909 = new_n18626_ | new_n18627_;
  assign new_n18629_ = pi028 & new_n18326_;
  assign new_n18630_ = ~pi028 & lo0910;
  assign li0910 = new_n18629_ | new_n18630_;
  assign new_n18632_ = pi041 & new_n18326_;
  assign new_n18633_ = ~pi041 & lo0911;
  assign li0911 = new_n18632_ | new_n18633_;
  assign new_n18635_ = pi025 & new_n18326_;
  assign new_n18636_ = ~pi025 & lo0912;
  assign li0912 = new_n18635_ | new_n18636_;
  assign new_n18638_ = pi017 & new_n18326_;
  assign new_n18639_ = ~pi017 & lo0913;
  assign li0913 = new_n18638_ | new_n18639_;
  assign new_n18641_ = ~lo0280 & new_n17052_;
  assign new_n18642_ = lo0280 & ~new_n17052_;
  assign li0914 = new_n18641_ | new_n18642_;
  assign new_n18644_ = pi019 & new_n18326_;
  assign new_n18645_ = ~pi019 & lo0915;
  assign li0915 = new_n18644_ | new_n18645_;
  assign new_n18647_ = pi034 & new_n18326_;
  assign new_n18648_ = ~pi034 & lo0916;
  assign li0916 = new_n18647_ | new_n18648_;
  assign new_n18650_ = pi023 & new_n18326_;
  assign new_n18651_ = ~pi023 & lo0917;
  assign li0917 = new_n18650_ | new_n18651_;
  assign new_n18653_ = pi015 & new_n18326_;
  assign new_n18654_ = ~pi015 & lo0918;
  assign li0918 = new_n18653_ | new_n18654_;
  assign new_n18656_ = pi013 & new_n18326_;
  assign new_n18657_ = ~pi013 & lo0919;
  assign li0919 = new_n18656_ | new_n18657_;
  assign new_n18659_ = pi004 & lo0920;
  assign new_n18660_ = pi050 & ~lo0920;
  assign li0920 = new_n18659_ | new_n18660_;
  assign new_n18662_ = pi004 & lo0921;
  assign new_n18663_ = pi051 & ~lo0921;
  assign li0921 = new_n18662_ | new_n18663_;
  assign new_n18665_ = pi004 & lo0922;
  assign new_n18666_ = pi063 & ~lo0922;
  assign li0922 = new_n18665_ | new_n18666_;
  assign new_n18668_ = pi004 & lo0923;
  assign new_n18669_ = pi065 & ~lo0923;
  assign li0923 = new_n18668_ | new_n18669_;
  assign new_n18671_ = ~lo0311 & new_n15353_;
  assign li0924 = ~lo0301 & new_n18671_;
  assign new_n18673_ = pi004 & lo0925;
  assign new_n18674_ = pi066 & ~lo0925;
  assign li0925 = new_n18673_ | new_n18674_;
  assign new_n18676_ = pi004 & lo0926;
  assign new_n18677_ = pi068 & ~lo0926;
  assign li0926 = new_n18676_ | new_n18677_;
  assign new_n18679_ = pi004 & lo0927;
  assign new_n18680_ = pi056 & ~lo0927;
  assign li0927 = new_n18679_ | new_n18680_;
  assign new_n18682_ = pi004 & lo0928;
  assign new_n18683_ = pi047 & ~lo0928;
  assign li0928 = new_n18682_ | new_n18683_;
  assign new_n18685_ = pi004 & lo0929;
  assign new_n18686_ = pi055 & ~lo0929;
  assign li0929 = new_n18685_ | new_n18686_;
  assign new_n18688_ = pi004 & lo0930;
  assign new_n18689_ = pi045 & ~lo0930;
  assign li0930 = new_n18688_ | new_n18689_;
  assign new_n18691_ = pi004 & lo0931;
  assign new_n18692_ = pi061 & ~lo0931;
  assign li0931 = new_n18691_ | new_n18692_;
  assign new_n18694_ = pi004 & lo0932;
  assign new_n18695_ = pi053 & ~lo0932;
  assign li0932 = new_n18694_ | new_n18695_;
  assign new_n18697_ = pi004 & lo0933;
  assign new_n18698_ = pi048 & ~lo0933;
  assign li0933 = new_n18697_ | new_n18698_;
  assign new_n18700_ = pi004 & lo0934;
  assign new_n18701_ = pi058 & ~lo0934;
  assign li0934 = new_n18700_ | new_n18701_;
  assign new_n18703_ = pi004 & lo0935;
  assign new_n18704_ = pi052 & ~lo0935;
  assign li0935 = new_n18703_ | new_n18704_;
  assign new_n18706_ = pi004 & lo0936;
  assign new_n18707_ = pi060 & ~lo0936;
  assign li0936 = new_n18706_ | new_n18707_;
  assign new_n18709_ = pi004 & lo0937;
  assign new_n18710_ = pi059 & ~lo0937;
  assign li0937 = new_n18709_ | new_n18710_;
  assign new_n18712_ = pi004 & lo0938;
  assign new_n18713_ = pi046 & ~lo0938;
  assign li0938 = new_n18712_ | new_n18713_;
  assign new_n18715_ = pi004 & lo0939;
  assign new_n18716_ = pi057 & ~lo0939;
  assign li0939 = new_n18715_ | new_n18716_;
  assign new_n18718_ = pi004 & lo0940;
  assign new_n18719_ = pi049 & ~lo0940;
  assign li0940 = new_n18718_ | new_n18719_;
  assign new_n18721_ = pi004 & lo0941;
  assign new_n18722_ = pi064 & ~lo0941;
  assign li0941 = new_n18721_ | new_n18722_;
  assign new_n18724_ = pi004 & lo0942;
  assign new_n18725_ = pi067 & ~lo0942;
  assign li0942 = new_n18724_ | new_n18725_;
  assign new_n18727_ = pi004 & lo0943;
  assign new_n18728_ = pi062 & ~lo0943;
  assign li0943 = new_n18727_ | new_n18728_;
  assign new_n18730_ = pi004 & lo0944;
  assign new_n18731_ = pi054 & ~lo0944;
  assign li0944 = new_n18730_ | new_n18731_;
  assign li0945 = new_n4454_ | new_n4466_;
  assign new_n18734_ = lo0782 & ~new_n18618_;
  assign new_n18735_ = ~lo0782 & lo0947;
  assign li0947 = new_n18734_ | new_n18735_;
  assign new_n18737_ = ~lo0266 & new_n17051_;
  assign new_n18738_ = lo0266 & ~new_n17051_;
  assign li0948 = new_n18737_ | new_n18738_;
  assign new_n18740_ = lo0949 & ~lo0954;
  assign new_n18741_ = lo0313 & ~lo0949;
  assign li0949 = new_n18740_ | new_n18741_;
  assign new_n18743_ = pi003 & lo0957;
  assign li0957 = lo0031 | new_n18743_;
  assign new_n18745_ = ~lo0278 & lo0279;
  assign new_n18746_ = lo0278 & ~lo0279;
  assign li0958 = new_n18745_ | new_n18746_;
  assign li0960 = ~lo0782 & lo0960;
  assign li0961 = ~lo0230 & lo0961;
  assign li0963 = ~lo0782 & lo0963;
  assign li0967 = ~lo0230 & lo0967;
  assign li0969 = ~lo0230 & lo0969;
  assign li0970 = ~lo0782 & lo0970;
  assign li0971 = ~lo0230 & lo0971;
  assign li0972 = ~lo0782 & lo0972;
  assign li0974 = ~lo0230 & lo0974;
  assign li0975 = ~lo0782 & lo0975;
  assign li0977 = ~lo0230 & lo0977;
  assign li0978 = ~lo0782 & lo0978;
  assign li0979 = lo0598 | lo0615;
  assign li0984 = lo0604 | lo0624;
  assign li0998 = 1'b0;
  assign li1001 = 1'b0;
  assign li1008 = 1'b0;
  assign li1023 = 1'b0;
  assign li0954 = ~lo0954;
  assign li0976 = ~lo0278;
  assign po000 = lo0668;
  assign po001 = lo0672;
  assign po002 = lo0664;
  assign po003 = lo0667;
  assign po004 = lo0676;
  assign po005 = lo0673;
  assign po006 = lo0675;
  assign po007 = lo0666;
  assign po008 = lo0679;
  assign po009 = lo0674;
  assign po010 = lo0663;
  assign po011 = lo0670;
  assign po012 = lo0677;
  assign po013 = lo0682;
  assign po014 = lo0671;
  assign po015 = lo0678;
  assign po016 = lo0718;
  assign po017 = lo0707;
  assign po018 = lo0708;
  assign po019 = lo0713;
  assign po020 = lo0711;
  assign po021 = lo0716;
  assign po022 = lo0733;
  assign po023 = lo0712;
  assign po024 = lo0689;
  assign po025 = lo0717;
  assign po026 = lo0692;
  assign po027 = lo0719;
  assign po028 = lo0722;
  assign po029 = lo0714;
  assign po030 = lo0720;
  assign po031 = lo0685;
  assign po032 = lo0837;
  assign po033 = lo0850;
  assign po034 = lo0872;
  assign po035 = lo0871;
  assign po036 = lo0881;
  assign po037 = lo0866;
  assign po038 = lo0876;
  assign po039 = lo0873;
  assign po040 = lo0874;
  assign po041 = lo0859;
  assign po042 = lo0855;
  assign po043 = lo0852;
  assign po044 = lo0870;
  assign po045 = lo0848;
  assign po046 = lo0865;
  assign po047 = lo0856;
  assign po048 = lo0853;
  assign po049 = lo0847;
  assign po050 = lo0857;
  assign po051 = lo0854;
  assign po052 = lo0858;
  assign po053 = lo0845;
  assign po054 = lo0838;
  assign po055 = lo0842;
  assign po056 = lo0843;
  assign po057 = lo0839;
  assign po058 = lo0844;
  assign po059 = lo0868;
  assign po060 = lo0851;
  assign po061 = lo0867;
  assign po062 = lo0880;
  assign po063 = lo0860;
  assign po064 = lo1024;
  assign po065 = lo1028;
  assign po066 = lo1009;
  assign po067 = lo1014;
  assign po068 = lo1019;
  assign po069 = lo0999;
  assign po070 = lo0990;
  assign po071 = lo1006;
  assign po072 = lo0987;
  assign po073 = lo1010;
  assign po074 = lo1015;
  assign po075 = lo1004;
  assign po076 = lo1021;
  assign po077 = lo1012;
  assign po078 = lo1011;
  assign po079 = lo1018;
  assign po080 = lo1003;
  assign po081 = lo1026;
  assign po082 = lo0997;
  assign po083 = lo0991;
  assign po084 = lo1007;
  assign po085 = lo1005;
  assign po086 = lo1002;
  assign po087 = lo1013;
  assign po088 = lo1025;
  assign po089 = lo1016;
  assign po090 = lo0994;
  assign po091 = lo1017;
  assign po092 = lo0996;
  assign po093 = lo1020;
  assign po094 = lo1000;
  assign po095 = lo0992;
  assign po096 = lo0031;
  assign po097 = lo0080;
  assign po098 = lo0893;
  assign po099 = lo0467;
  assign po100 = lo0078;
  assign po101 = lo0112;
  assign po102 = lo0013;
  assign po103 = lo0025;
  assign po104 = lo0226;
  assign po105 = lo0127;
  assign po106 = lo0822;
  assign po107 = lo0808;
  assign po108 = lo0227;
  assign po109 = lo0477;
  assign po110 = lo0834;
  assign po111 = lo0229;
  assign po112 = lo0012;
  assign po113 = lo0011;
  assign po114 = lo0010;
  assign po115 = lo0009;
  assign po116 = lo0008;
  assign po117 = lo0007;
  assign po118 = lo0006;
  assign po119 = lo0005;
  assign po120 = lo0004;
  assign po121 = lo0003;
  assign po122 = lo0000;
  assign po123 = lo0002;
  assign po124 = lo0001;
  assign po125 = lo0310;
  assign po126 = lo0302;
  assign po127 = lo0475;
  assign po128 = lo0474;
  assign po129 = lo0466;
  assign po130 = lo0473;
  assign po131 = lo0471;
  assign po132 = lo0472;
  assign po133 = lo0470;
  assign po134 = lo0469;
  assign po135 = lo0465;
  assign po136 = lo1022;
  assign po137 = lo1027;
  assign po138 = lo0989;
  assign po139 = lo0988;
  assign po140 = lo0028;
  assign po141 = lo0027;
  assign po142 = lo0026;
  assign po143 = lo0029;
  assign po144 = lo0015;
  assign po145 = lo0014;
  assign po146 = lo0021;
  assign po147 = lo0020;
  assign po148 = lo0019;
  assign po149 = lo0018;
  assign po150 = lo0017;
  assign po151 = lo0016;
  assign li0022 = lo0023;
  assign li0023 = li0013;
  assign li0030 = lo0037;
  assign li0105 = lo0117;
  assign li0123 = li0122;
  assign li0128 = lo0131;
  assign li0229 = lo0232;
  assign li0231 = lo0236;
  assign li0479 = lo0583;
  assign li0834 = lo0893;
  assign li0897 = lo0067;
  assign li0952 = pi045;
  assign li0953 = pi045;
  assign li0955 = lo0965;
  assign li0956 = pi045;
  assign li0959 = lo0985;
  assign li0962 = lo1008;
  assign li0964 = lo1023;
  assign li0965 = lo0998;
  assign li0966 = lo1001;
  assign li0968 = pi046;
  assign li0973 = pi046;
  assign li0980 = pi046;
  assign li0981 = lo1058;
  assign li0983 = lo0299;
  assign li0985 = lo1069;
  assign li0986 = lo1046;
  assign li0987 = lo0915;
  assign li0988 = lo0825;
  assign li0989 = lo0826;
  assign li0990 = lo0913;
  assign li0991 = lo0894;
  assign li0992 = lo0905;
  assign li0993 = pi006;
  assign li0994 = lo0890;
  assign li0995 = pi005;
  assign li0996 = lo0906;
  assign li0997 = lo0896;
  assign li0999 = lo0909;
  assign li1000 = lo0911;
  assign li1002 = lo0908;
  assign li1003 = lo0891;
  assign li1004 = lo0902;
  assign li1005 = lo0903;
  assign li1006 = lo0883;
  assign li1007 = lo0888;
  assign li1009 = lo0919;
  assign li1010 = lo0886;
  assign li1011 = lo0912;
  assign li1012 = lo0895;
  assign li1013 = lo0916;
  assign li1014 = lo0889;
  assign li1015 = lo0900;
  assign li1016 = lo0885;
  assign li1017 = lo0904;
  assign li1018 = lo0899;
  assign li1019 = lo0918;
  assign li1020 = lo0898;
  assign li1021 = lo0917;
  assign li1022 = lo0827;
  assign li1024 = lo0887;
  assign li1025 = lo0884;
  assign li1026 = lo0910;
  assign li1027 = lo0828;
  assign li1028 = lo0892;
  assign li1029 = pi098;
  assign li1030 = pi083;
  assign li1031 = pi081;
  assign li1032 = pi049;
  assign li1033 = pi088;
  assign li1034 = pi089;
  assign li1035 = lo0863;
  assign li1036 = pi114;
  assign li1037 = pi096;
  assign li1038 = pi082;
  assign li1039 = pi103;
  assign li1040 = pi048;
  assign li1041 = pi097;
  assign li1042 = pi076;
  assign li1043 = pi075;
  assign li1044 = pi009;
  assign li1045 = pi094;
  assign li1046 = lo0230;
  assign li1047 = pi080;
  assign li1048 = pi047;
  assign li1049 = pi092;
  assign li1050 = lo0849;
  assign li1051 = pi104;
  assign li1052 = pi093;
  assign li1053 = pi079;
  assign li1054 = pi048;
  assign li1055 = pi047;
  assign li1056 = pi086;
  assign li1057 = pi102;
  assign li1058 = pi010;
  assign li1059 = pi085;
  assign li1060 = pi048;
  assign li1061 = pi090;
  assign li1062 = pi113;
  assign li1063 = pi087;
  assign li1064 = pi084;
  assign li1065 = pi112;
  assign li1066 = pi078;
  assign li1067 = lo0840;
  assign li1068 = pi100;
  assign li1069 = lo0127;
  assign li1070 = pi106;
  assign li1071 = lo0864;
  assign li1072 = pi101;
  assign li1073 = pi099;
  assign li1074 = pi091;
  assign li1075 = pi105;
  assign li1076 = pi008;
  assign li1077 = pi049;
  assign li1078 = pi077;
  assign li1079 = pi047;
  assign li1080 = pi111;
  assign li1081 = pi095;
  assign li1082 = pi049;
  always @ (posedge clock) begin
    lo0000 <= li0000;
    lo0001 <= li0001;
    lo0002 <= li0002;
    lo0003 <= li0003;
    lo0004 <= li0004;
    lo0005 <= li0005;
    lo0006 <= li0006;
    lo0007 <= li0007;
    lo0008 <= li0008;
    lo0009 <= li0009;
    lo0010 <= li0010;
    lo0011 <= li0011;
    lo0012 <= li0012;
    lo0013 <= li0013;
    lo0014 <= li0014;
    lo0015 <= li0015;
    lo0016 <= li0016;
    lo0017 <= li0017;
    lo0018 <= li0018;
    lo0019 <= li0019;
    lo0020 <= li0020;
    lo0021 <= li0021;
    lo0022 <= li0022;
    lo0023 <= li0023;
    lo0024 <= li0024;
    lo0025 <= li0025;
    lo0026 <= li0026;
    lo0027 <= li0027;
    lo0028 <= li0028;
    lo0029 <= li0029;
    lo0030 <= li0030;
    lo0031 <= li0031;
    lo0032 <= li0032;
    lo0033 <= li0033;
    lo0034 <= li0034;
    lo0035 <= li0035;
    lo0036 <= li0036;
    lo0037 <= li0037;
    lo0038 <= li0038;
    lo0039 <= li0039;
    lo0040 <= li0040;
    lo0041 <= li0041;
    lo0042 <= li0042;
    lo0043 <= li0043;
    lo0044 <= li0044;
    lo0045 <= li0045;
    lo0046 <= li0046;
    lo0047 <= li0047;
    lo0048 <= li0048;
    lo0049 <= li0049;
    lo0050 <= li0050;
    lo0051 <= li0051;
    lo0052 <= li0052;
    lo0053 <= li0053;
    lo0054 <= li0054;
    lo0055 <= li0055;
    lo0056 <= li0056;
    lo0057 <= li0057;
    lo0058 <= li0058;
    lo0059 <= li0059;
    lo0060 <= li0060;
    lo0061 <= li0061;
    lo0062 <= li0062;
    lo0063 <= li0063;
    lo0064 <= li0064;
    lo0065 <= li0065;
    lo0066 <= li0066;
    lo0067 <= li0067;
    lo0068 <= li0068;
    lo0069 <= li0069;
    lo0070 <= li0070;
    lo0071 <= li0071;
    lo0072 <= li0072;
    lo0073 <= li0073;
    lo0074 <= li0074;
    lo0075 <= li0075;
    lo0076 <= li0076;
    lo0077 <= li0077;
    lo0078 <= li0078;
    lo0079 <= li0079;
    lo0080 <= li0080;
    lo0081 <= li0081;
    lo0082 <= li0082;
    lo0083 <= li0083;
    lo0084 <= li0084;
    lo0085 <= li0085;
    lo0086 <= li0086;
    lo0087 <= li0087;
    lo0088 <= li0088;
    lo0089 <= li0089;
    lo0090 <= li0090;
    lo0091 <= li0091;
    lo0092 <= li0092;
    lo0093 <= li0093;
    lo0094 <= li0094;
    lo0095 <= li0095;
    lo0096 <= li0096;
    lo0097 <= li0097;
    lo0098 <= li0098;
    lo0099 <= li0099;
    lo0100 <= li0100;
    lo0101 <= li0101;
    lo0102 <= li0102;
    lo0103 <= li0103;
    lo0104 <= li0104;
    lo0105 <= li0105;
    lo0106 <= li0106;
    lo0107 <= li0107;
    lo0108 <= li0108;
    lo0109 <= li0109;
    lo0110 <= li0110;
    lo0111 <= li0111;
    lo0112 <= li0112;
    lo0113 <= li0113;
    lo0114 <= li0114;
    lo0115 <= li0115;
    lo0116 <= li0116;
    lo0117 <= li0117;
    lo0118 <= li0118;
    lo0119 <= li0119;
    lo0120 <= li0120;
    lo0121 <= li0121;
    lo0122 <= li0122;
    lo0123 <= li0123;
    lo0124 <= li0124;
    lo0125 <= li0125;
    lo0126 <= li0126;
    lo0127 <= li0127;
    lo0128 <= li0128;
    lo0129 <= li0129;
    lo0130 <= li0130;
    lo0131 <= li0131;
    lo0132 <= li0132;
    lo0133 <= li0133;
    lo0134 <= li0134;
    lo0135 <= li0135;
    lo0136 <= li0136;
    lo0137 <= li0137;
    lo0138 <= li0138;
    lo0139 <= li0139;
    lo0140 <= li0140;
    lo0141 <= li0141;
    lo0142 <= li0142;
    lo0143 <= li0143;
    lo0144 <= li0144;
    lo0145 <= li0145;
    lo0146 <= li0146;
    lo0147 <= li0147;
    lo0148 <= li0148;
    lo0149 <= li0149;
    lo0150 <= li0150;
    lo0151 <= li0151;
    lo0152 <= li0152;
    lo0153 <= li0153;
    lo0154 <= li0154;
    lo0155 <= li0155;
    lo0156 <= li0156;
    lo0157 <= li0157;
    lo0158 <= li0158;
    lo0159 <= li0159;
    lo0160 <= li0160;
    lo0161 <= li0161;
    lo0162 <= li0162;
    lo0163 <= li0163;
    lo0164 <= li0164;
    lo0165 <= li0165;
    lo0166 <= li0166;
    lo0167 <= li0167;
    lo0168 <= li0168;
    lo0169 <= li0169;
    lo0170 <= li0170;
    lo0171 <= li0171;
    lo0172 <= li0172;
    lo0173 <= li0173;
    lo0174 <= li0174;
    lo0175 <= li0175;
    lo0176 <= li0176;
    lo0177 <= li0177;
    lo0178 <= li0178;
    lo0179 <= li0179;
    lo0180 <= li0180;
    lo0181 <= li0181;
    lo0182 <= li0182;
    lo0183 <= li0183;
    lo0184 <= li0184;
    lo0185 <= li0185;
    lo0186 <= li0186;
    lo0187 <= li0187;
    lo0188 <= li0188;
    lo0189 <= li0189;
    lo0190 <= li0190;
    lo0191 <= li0191;
    lo0192 <= li0192;
    lo0193 <= li0193;
    lo0194 <= li0194;
    lo0195 <= li0195;
    lo0196 <= li0196;
    lo0197 <= li0197;
    lo0198 <= li0198;
    lo0199 <= li0199;
    lo0200 <= li0200;
    lo0201 <= li0201;
    lo0202 <= li0202;
    lo0203 <= li0203;
    lo0204 <= li0204;
    lo0205 <= li0205;
    lo0206 <= li0206;
    lo0207 <= li0207;
    lo0208 <= li0208;
    lo0209 <= li0209;
    lo0210 <= li0210;
    lo0211 <= li0211;
    lo0212 <= li0212;
    lo0213 <= li0213;
    lo0214 <= li0214;
    lo0215 <= li0215;
    lo0216 <= li0216;
    lo0217 <= li0217;
    lo0218 <= li0218;
    lo0219 <= li0219;
    lo0220 <= li0220;
    lo0221 <= li0221;
    lo0222 <= li0222;
    lo0223 <= li0223;
    lo0224 <= li0224;
    lo0225 <= li0225;
    lo0226 <= li0226;
    lo0227 <= li0227;
    lo0228 <= li0228;
    lo0229 <= li0229;
    lo0230 <= li0230;
    lo0231 <= li0231;
    lo0232 <= li0232;
    lo0233 <= li0233;
    lo0234 <= li0234;
    lo0235 <= li0235;
    lo0236 <= li0236;
    lo0237 <= li0237;
    lo0238 <= li0238;
    lo0239 <= li0239;
    lo0240 <= li0240;
    lo0241 <= li0241;
    lo0242 <= li0242;
    lo0243 <= li0243;
    lo0244 <= li0244;
    lo0245 <= li0245;
    lo0246 <= li0246;
    lo0247 <= li0247;
    lo0248 <= li0248;
    lo0249 <= li0249;
    lo0250 <= li0250;
    lo0251 <= li0251;
    lo0252 <= li0252;
    lo0253 <= li0253;
    lo0254 <= li0254;
    lo0255 <= li0255;
    lo0256 <= li0256;
    lo0257 <= li0257;
    lo0258 <= li0258;
    lo0259 <= li0259;
    lo0260 <= li0260;
    lo0261 <= li0261;
    lo0262 <= li0262;
    lo0263 <= li0263;
    lo0264 <= li0264;
    lo0265 <= li0265;
    lo0266 <= li0266;
    lo0267 <= li0267;
    lo0268 <= li0268;
    lo0269 <= li0269;
    lo0270 <= li0270;
    lo0271 <= li0271;
    lo0272 <= li0272;
    lo0273 <= li0273;
    lo0274 <= li0274;
    lo0275 <= li0275;
    lo0276 <= li0276;
    lo0277 <= li0277;
    lo0278 <= li0278;
    lo0279 <= li0279;
    lo0280 <= li0280;
    lo0281 <= li0281;
    lo0282 <= li0282;
    lo0283 <= li0283;
    lo0284 <= li0284;
    lo0285 <= li0285;
    lo0286 <= li0286;
    lo0287 <= li0287;
    lo0288 <= li0288;
    lo0289 <= li0289;
    lo0290 <= li0290;
    lo0291 <= li0291;
    lo0292 <= li0292;
    lo0293 <= li0293;
    lo0294 <= li0294;
    lo0295 <= li0295;
    lo0296 <= li0296;
    lo0297 <= li0297;
    lo0298 <= li0298;
    lo0299 <= li0299;
    lo0300 <= li0300;
    lo0301 <= li0301;
    lo0302 <= li0302;
    lo0303 <= li0303;
    lo0304 <= li0304;
    lo0305 <= li0305;
    lo0306 <= li0306;
    lo0307 <= li0307;
    lo0308 <= li0308;
    lo0309 <= li0309;
    lo0310 <= li0310;
    lo0311 <= li0311;
    lo0312 <= li0312;
    lo0313 <= li0313;
    lo0314 <= li0314;
    lo0315 <= li0315;
    lo0316 <= li0316;
    lo0317 <= li0317;
    lo0318 <= li0318;
    lo0319 <= li0319;
    lo0320 <= li0320;
    lo0321 <= li0321;
    lo0322 <= li0322;
    lo0323 <= li0323;
    lo0324 <= li0324;
    lo0325 <= li0325;
    lo0326 <= li0326;
    lo0327 <= li0327;
    lo0328 <= li0328;
    lo0329 <= li0329;
    lo0330 <= li0330;
    lo0331 <= li0331;
    lo0332 <= li0332;
    lo0333 <= li0333;
    lo0334 <= li0334;
    lo0335 <= li0335;
    lo0336 <= li0336;
    lo0337 <= li0337;
    lo0338 <= li0338;
    lo0339 <= li0339;
    lo0340 <= li0340;
    lo0341 <= li0341;
    lo0342 <= li0342;
    lo0343 <= li0343;
    lo0344 <= li0344;
    lo0345 <= li0345;
    lo0346 <= li0346;
    lo0347 <= li0347;
    lo0348 <= li0348;
    lo0349 <= li0349;
    lo0350 <= li0350;
    lo0351 <= li0351;
    lo0352 <= li0352;
    lo0353 <= li0353;
    lo0354 <= li0354;
    lo0355 <= li0355;
    lo0356 <= li0356;
    lo0357 <= li0357;
    lo0358 <= li0358;
    lo0359 <= li0359;
    lo0360 <= li0360;
    lo0361 <= li0361;
    lo0362 <= li0362;
    lo0363 <= li0363;
    lo0364 <= li0364;
    lo0365 <= li0365;
    lo0366 <= li0366;
    lo0367 <= li0367;
    lo0368 <= li0368;
    lo0369 <= li0369;
    lo0370 <= li0370;
    lo0371 <= li0371;
    lo0372 <= li0372;
    lo0373 <= li0373;
    lo0374 <= li0374;
    lo0375 <= li0375;
    lo0376 <= li0376;
    lo0377 <= li0377;
    lo0378 <= li0378;
    lo0379 <= li0379;
    lo0380 <= li0380;
    lo0381 <= li0381;
    lo0382 <= li0382;
    lo0383 <= li0383;
    lo0384 <= li0384;
    lo0385 <= li0385;
    lo0386 <= li0386;
    lo0387 <= li0387;
    lo0388 <= li0388;
    lo0389 <= li0389;
    lo0390 <= li0390;
    lo0391 <= li0391;
    lo0392 <= li0392;
    lo0393 <= li0393;
    lo0394 <= li0394;
    lo0395 <= li0395;
    lo0396 <= li0396;
    lo0397 <= li0397;
    lo0398 <= li0398;
    lo0399 <= li0399;
    lo0400 <= li0400;
    lo0401 <= li0401;
    lo0402 <= li0402;
    lo0403 <= li0403;
    lo0404 <= li0404;
    lo0405 <= li0405;
    lo0406 <= li0406;
    lo0407 <= li0407;
    lo0408 <= li0408;
    lo0409 <= li0409;
    lo0410 <= li0410;
    lo0411 <= li0411;
    lo0412 <= li0412;
    lo0413 <= li0413;
    lo0414 <= li0414;
    lo0415 <= li0415;
    lo0416 <= li0416;
    lo0417 <= li0417;
    lo0418 <= li0418;
    lo0419 <= li0419;
    lo0420 <= li0420;
    lo0421 <= li0421;
    lo0422 <= li0422;
    lo0423 <= li0423;
    lo0424 <= li0424;
    lo0425 <= li0425;
    lo0426 <= li0426;
    lo0427 <= li0427;
    lo0428 <= li0428;
    lo0429 <= li0429;
    lo0430 <= li0430;
    lo0431 <= li0431;
    lo0432 <= li0432;
    lo0433 <= li0433;
    lo0434 <= li0434;
    lo0435 <= li0435;
    lo0436 <= li0436;
    lo0437 <= li0437;
    lo0438 <= li0438;
    lo0439 <= li0439;
    lo0440 <= li0440;
    lo0441 <= li0441;
    lo0442 <= li0442;
    lo0443 <= li0443;
    lo0444 <= li0444;
    lo0445 <= li0445;
    lo0446 <= li0446;
    lo0447 <= li0447;
    lo0448 <= li0448;
    lo0449 <= li0449;
    lo0450 <= li0450;
    lo0451 <= li0451;
    lo0452 <= li0452;
    lo0453 <= li0453;
    lo0454 <= li0454;
    lo0455 <= li0455;
    lo0456 <= li0456;
    lo0457 <= li0457;
    lo0458 <= li0458;
    lo0459 <= li0459;
    lo0460 <= li0460;
    lo0461 <= li0461;
    lo0462 <= li0462;
    lo0463 <= li0463;
    lo0464 <= li0464;
    lo0465 <= li0465;
    lo0466 <= li0466;
    lo0467 <= li0467;
    lo0468 <= li0468;
    lo0469 <= li0469;
    lo0470 <= li0470;
    lo0471 <= li0471;
    lo0472 <= li0472;
    lo0473 <= li0473;
    lo0474 <= li0474;
    lo0475 <= li0475;
    lo0476 <= li0476;
    lo0477 <= li0477;
    lo0478 <= li0478;
    lo0479 <= li0479;
    lo0480 <= li0480;
    lo0481 <= li0481;
    lo0482 <= li0482;
    lo0483 <= li0483;
    lo0484 <= li0484;
    lo0485 <= li0485;
    lo0486 <= li0486;
    lo0487 <= li0487;
    lo0488 <= li0488;
    lo0489 <= li0489;
    lo0490 <= li0490;
    lo0491 <= li0491;
    lo0492 <= li0492;
    lo0493 <= li0493;
    lo0494 <= li0494;
    lo0495 <= li0495;
    lo0496 <= li0496;
    lo0497 <= li0497;
    lo0498 <= li0498;
    lo0499 <= li0499;
    lo0500 <= li0500;
    lo0501 <= li0501;
    lo0502 <= li0502;
    lo0503 <= li0503;
    lo0504 <= li0504;
    lo0505 <= li0505;
    lo0506 <= li0506;
    lo0507 <= li0507;
    lo0508 <= li0508;
    lo0509 <= li0509;
    lo0510 <= li0510;
    lo0511 <= li0511;
    lo0512 <= li0512;
    lo0513 <= li0513;
    lo0514 <= li0514;
    lo0515 <= li0515;
    lo0516 <= li0516;
    lo0517 <= li0517;
    lo0518 <= li0518;
    lo0519 <= li0519;
    lo0520 <= li0520;
    lo0521 <= li0521;
    lo0522 <= li0522;
    lo0523 <= li0523;
    lo0524 <= li0524;
    lo0525 <= li0525;
    lo0526 <= li0526;
    lo0527 <= li0527;
    lo0528 <= li0528;
    lo0529 <= li0529;
    lo0530 <= li0530;
    lo0531 <= li0531;
    lo0532 <= li0532;
    lo0533 <= li0533;
    lo0534 <= li0534;
    lo0535 <= li0535;
    lo0536 <= li0536;
    lo0537 <= li0537;
    lo0538 <= li0538;
    lo0539 <= li0539;
    lo0540 <= li0540;
    lo0541 <= li0541;
    lo0542 <= li0542;
    lo0543 <= li0543;
    lo0544 <= li0544;
    lo0545 <= li0545;
    lo0546 <= li0546;
    lo0547 <= li0547;
    lo0548 <= li0548;
    lo0549 <= li0549;
    lo0550 <= li0550;
    lo0551 <= li0551;
    lo0552 <= li0552;
    lo0553 <= li0553;
    lo0554 <= li0554;
    lo0555 <= li0555;
    lo0556 <= li0556;
    lo0557 <= li0557;
    lo0558 <= li0558;
    lo0559 <= li0559;
    lo0560 <= li0560;
    lo0561 <= li0561;
    lo0562 <= li0562;
    lo0563 <= li0563;
    lo0564 <= li0564;
    lo0565 <= li0565;
    lo0566 <= li0566;
    lo0567 <= li0567;
    lo0568 <= li0568;
    lo0569 <= li0569;
    lo0570 <= li0570;
    lo0571 <= li0571;
    lo0572 <= li0572;
    lo0573 <= li0573;
    lo0574 <= li0574;
    lo0575 <= li0575;
    lo0576 <= li0576;
    lo0577 <= li0577;
    lo0578 <= li0578;
    lo0579 <= li0579;
    lo0580 <= li0580;
    lo0581 <= li0581;
    lo0582 <= li0582;
    lo0583 <= li0583;
    lo0584 <= li0584;
    lo0585 <= li0585;
    lo0586 <= li0586;
    lo0587 <= li0587;
    lo0588 <= li0588;
    lo0589 <= li0589;
    lo0590 <= li0590;
    lo0591 <= li0591;
    lo0592 <= li0592;
    lo0593 <= li0593;
    lo0594 <= li0594;
    lo0595 <= li0595;
    lo0596 <= li0596;
    lo0597 <= li0597;
    lo0598 <= li0598;
    lo0599 <= li0599;
    lo0600 <= li0600;
    lo0601 <= li0601;
    lo0602 <= li0602;
    lo0603 <= li0603;
    lo0604 <= li0604;
    lo0605 <= li0605;
    lo0606 <= li0606;
    lo0607 <= li0607;
    lo0608 <= li0608;
    lo0609 <= li0609;
    lo0610 <= li0610;
    lo0611 <= li0611;
    lo0612 <= li0612;
    lo0613 <= li0613;
    lo0614 <= li0614;
    lo0615 <= li0615;
    lo0616 <= li0616;
    lo0617 <= li0617;
    lo0618 <= li0618;
    lo0619 <= li0619;
    lo0620 <= li0620;
    lo0621 <= li0621;
    lo0622 <= li0622;
    lo0623 <= li0623;
    lo0624 <= li0624;
    lo0625 <= li0625;
    lo0626 <= li0626;
    lo0627 <= li0627;
    lo0628 <= li0628;
    lo0629 <= li0629;
    lo0630 <= li0630;
    lo0631 <= li0631;
    lo0632 <= li0632;
    lo0633 <= li0633;
    lo0634 <= li0634;
    lo0635 <= li0635;
    lo0636 <= li0636;
    lo0637 <= li0637;
    lo0638 <= li0638;
    lo0639 <= li0639;
    lo0640 <= li0640;
    lo0641 <= li0641;
    lo0642 <= li0642;
    lo0643 <= li0643;
    lo0644 <= li0644;
    lo0645 <= li0645;
    lo0646 <= li0646;
    lo0647 <= li0647;
    lo0648 <= li0648;
    lo0649 <= li0649;
    lo0650 <= li0650;
    lo0651 <= li0651;
    lo0652 <= li0652;
    lo0653 <= li0653;
    lo0654 <= li0654;
    lo0655 <= li0655;
    lo0656 <= li0656;
    lo0657 <= li0657;
    lo0658 <= li0658;
    lo0659 <= li0659;
    lo0660 <= li0660;
    lo0661 <= li0661;
    lo0662 <= li0662;
    lo0663 <= li0663;
    lo0664 <= li0664;
    lo0665 <= li0665;
    lo0666 <= li0666;
    lo0667 <= li0667;
    lo0668 <= li0668;
    lo0669 <= li0669;
    lo0670 <= li0670;
    lo0671 <= li0671;
    lo0672 <= li0672;
    lo0673 <= li0673;
    lo0674 <= li0674;
    lo0675 <= li0675;
    lo0676 <= li0676;
    lo0677 <= li0677;
    lo0678 <= li0678;
    lo0679 <= li0679;
    lo0680 <= li0680;
    lo0681 <= li0681;
    lo0682 <= li0682;
    lo0683 <= li0683;
    lo0684 <= li0684;
    lo0685 <= li0685;
    lo0686 <= li0686;
    lo0687 <= li0687;
    lo0688 <= li0688;
    lo0689 <= li0689;
    lo0690 <= li0690;
    lo0691 <= li0691;
    lo0692 <= li0692;
    lo0693 <= li0693;
    lo0694 <= li0694;
    lo0695 <= li0695;
    lo0696 <= li0696;
    lo0697 <= li0697;
    lo0698 <= li0698;
    lo0699 <= li0699;
    lo0700 <= li0700;
    lo0701 <= li0701;
    lo0702 <= li0702;
    lo0703 <= li0703;
    lo0704 <= li0704;
    lo0705 <= li0705;
    lo0706 <= li0706;
    lo0707 <= li0707;
    lo0708 <= li0708;
    lo0709 <= li0709;
    lo0710 <= li0710;
    lo0711 <= li0711;
    lo0712 <= li0712;
    lo0713 <= li0713;
    lo0714 <= li0714;
    lo0715 <= li0715;
    lo0716 <= li0716;
    lo0717 <= li0717;
    lo0718 <= li0718;
    lo0719 <= li0719;
    lo0720 <= li0720;
    lo0721 <= li0721;
    lo0722 <= li0722;
    lo0723 <= li0723;
    lo0724 <= li0724;
    lo0725 <= li0725;
    lo0726 <= li0726;
    lo0727 <= li0727;
    lo0728 <= li0728;
    lo0729 <= li0729;
    lo0730 <= li0730;
    lo0731 <= li0731;
    lo0732 <= li0732;
    lo0733 <= li0733;
    lo0734 <= li0734;
    lo0735 <= li0735;
    lo0736 <= li0736;
    lo0737 <= li0737;
    lo0738 <= li0738;
    lo0739 <= li0739;
    lo0740 <= li0740;
    lo0741 <= li0741;
    lo0742 <= li0742;
    lo0743 <= li0743;
    lo0744 <= li0744;
    lo0745 <= li0745;
    lo0746 <= li0746;
    lo0747 <= li0747;
    lo0748 <= li0748;
    lo0749 <= li0749;
    lo0750 <= li0750;
    lo0751 <= li0751;
    lo0752 <= li0752;
    lo0753 <= li0753;
    lo0754 <= li0754;
    lo0755 <= li0755;
    lo0756 <= li0756;
    lo0757 <= li0757;
    lo0758 <= li0758;
    lo0759 <= li0759;
    lo0760 <= li0760;
    lo0761 <= li0761;
    lo0762 <= li0762;
    lo0763 <= li0763;
    lo0764 <= li0764;
    lo0765 <= li0765;
    lo0766 <= li0766;
    lo0767 <= li0767;
    lo0768 <= li0768;
    lo0769 <= li0769;
    lo0770 <= li0770;
    lo0771 <= li0771;
    lo0772 <= li0772;
    lo0773 <= li0773;
    lo0774 <= li0774;
    lo0775 <= li0775;
    lo0776 <= li0776;
    lo0777 <= li0777;
    lo0778 <= li0778;
    lo0779 <= li0779;
    lo0780 <= li0780;
    lo0781 <= li0781;
    lo0782 <= li0782;
    lo0783 <= li0783;
    lo0784 <= li0784;
    lo0785 <= li0785;
    lo0786 <= li0786;
    lo0787 <= li0787;
    lo0788 <= li0788;
    lo0789 <= li0789;
    lo0790 <= li0790;
    lo0791 <= li0791;
    lo0792 <= li0792;
    lo0793 <= li0793;
    lo0794 <= li0794;
    lo0795 <= li0795;
    lo0796 <= li0796;
    lo0797 <= li0797;
    lo0798 <= li0798;
    lo0799 <= li0799;
    lo0800 <= li0800;
    lo0801 <= li0801;
    lo0802 <= li0802;
    lo0803 <= li0803;
    lo0804 <= li0804;
    lo0805 <= li0805;
    lo0806 <= li0806;
    lo0807 <= li0807;
    lo0808 <= li0808;
    lo0809 <= li0809;
    lo0810 <= li0810;
    lo0811 <= li0811;
    lo0812 <= li0812;
    lo0813 <= li0813;
    lo0814 <= li0814;
    lo0815 <= li0815;
    lo0816 <= li0816;
    lo0817 <= li0817;
    lo0818 <= li0818;
    lo0819 <= li0819;
    lo0820 <= li0820;
    lo0821 <= li0821;
    lo0822 <= li0822;
    lo0823 <= li0823;
    lo0824 <= li0824;
    lo0825 <= li0825;
    lo0826 <= li0826;
    lo0827 <= li0827;
    lo0828 <= li0828;
    lo0829 <= li0829;
    lo0830 <= li0830;
    lo0831 <= li0831;
    lo0832 <= li0832;
    lo0833 <= li0833;
    lo0834 <= li0834;
    lo0835 <= li0835;
    lo0836 <= li0836;
    lo0837 <= li0837;
    lo0838 <= li0838;
    lo0839 <= li0839;
    lo0840 <= li0840;
    lo0841 <= li0841;
    lo0842 <= li0842;
    lo0843 <= li0843;
    lo0844 <= li0844;
    lo0845 <= li0845;
    lo0846 <= li0846;
    lo0847 <= li0847;
    lo0848 <= li0848;
    lo0849 <= li0849;
    lo0850 <= li0850;
    lo0851 <= li0851;
    lo0852 <= li0852;
    lo0853 <= li0853;
    lo0854 <= li0854;
    lo0855 <= li0855;
    lo0856 <= li0856;
    lo0857 <= li0857;
    lo0858 <= li0858;
    lo0859 <= li0859;
    lo0860 <= li0860;
    lo0861 <= li0861;
    lo0862 <= li0862;
    lo0863 <= li0863;
    lo0864 <= li0864;
    lo0865 <= li0865;
    lo0866 <= li0866;
    lo0867 <= li0867;
    lo0868 <= li0868;
    lo0869 <= li0869;
    lo0870 <= li0870;
    lo0871 <= li0871;
    lo0872 <= li0872;
    lo0873 <= li0873;
    lo0874 <= li0874;
    lo0875 <= li0875;
    lo0876 <= li0876;
    lo0877 <= li0877;
    lo0878 <= li0878;
    lo0879 <= li0879;
    lo0880 <= li0880;
    lo0881 <= li0881;
    lo0882 <= li0882;
    lo0883 <= li0883;
    lo0884 <= li0884;
    lo0885 <= li0885;
    lo0886 <= li0886;
    lo0887 <= li0887;
    lo0888 <= li0888;
    lo0889 <= li0889;
    lo0890 <= li0890;
    lo0891 <= li0891;
    lo0892 <= li0892;
    lo0893 <= li0893;
    lo0894 <= li0894;
    lo0895 <= li0895;
    lo0896 <= li0896;
    lo0897 <= li0897;
    lo0898 <= li0898;
    lo0899 <= li0899;
    lo0900 <= li0900;
    lo0901 <= li0901;
    lo0902 <= li0902;
    lo0903 <= li0903;
    lo0904 <= li0904;
    lo0905 <= li0905;
    lo0906 <= li0906;
    lo0907 <= li0907;
    lo0908 <= li0908;
    lo0909 <= li0909;
    lo0910 <= li0910;
    lo0911 <= li0911;
    lo0912 <= li0912;
    lo0913 <= li0913;
    lo0914 <= li0914;
    lo0915 <= li0915;
    lo0916 <= li0916;
    lo0917 <= li0917;
    lo0918 <= li0918;
    lo0919 <= li0919;
    lo0920 <= li0920;
    lo0921 <= li0921;
    lo0922 <= li0922;
    lo0923 <= li0923;
    lo0924 <= li0924;
    lo0925 <= li0925;
    lo0926 <= li0926;
    lo0927 <= li0927;
    lo0928 <= li0928;
    lo0929 <= li0929;
    lo0930 <= li0930;
    lo0931 <= li0931;
    lo0932 <= li0932;
    lo0933 <= li0933;
    lo0934 <= li0934;
    lo0935 <= li0935;
    lo0936 <= li0936;
    lo0937 <= li0937;
    lo0938 <= li0938;
    lo0939 <= li0939;
    lo0940 <= li0940;
    lo0941 <= li0941;
    lo0942 <= li0942;
    lo0943 <= li0943;
    lo0944 <= li0944;
    lo0945 <= li0945;
    lo0946 <= li0946;
    lo0947 <= li0947;
    lo0948 <= li0948;
    lo0949 <= li0949;
    lo0950 <= li0950;
    lo0951 <= li0951;
    lo0952 <= li0952;
    lo0953 <= li0953;
    lo0954 <= li0954;
    lo0955 <= li0955;
    lo0956 <= li0956;
    lo0957 <= li0957;
    lo0958 <= li0958;
    lo0959 <= li0959;
    lo0960 <= li0960;
    lo0961 <= li0961;
    lo0962 <= li0962;
    lo0963 <= li0963;
    lo0964 <= li0964;
    lo0965 <= li0965;
    lo0966 <= li0966;
    lo0967 <= li0967;
    lo0968 <= li0968;
    lo0969 <= li0969;
    lo0970 <= li0970;
    lo0971 <= li0971;
    lo0972 <= li0972;
    lo0973 <= li0973;
    lo0974 <= li0974;
    lo0975 <= li0975;
    lo0976 <= li0976;
    lo0977 <= li0977;
    lo0978 <= li0978;
    lo0979 <= li0979;
    lo0980 <= li0980;
    lo0981 <= li0981;
    lo0982 <= li0982;
    lo0983 <= li0983;
    lo0984 <= li0984;
    lo0985 <= li0985;
    lo0986 <= li0986;
    lo0987 <= li0987;
    lo0988 <= li0988;
    lo0989 <= li0989;
    lo0990 <= li0990;
    lo0991 <= li0991;
    lo0992 <= li0992;
    lo0993 <= li0993;
    lo0994 <= li0994;
    lo0995 <= li0995;
    lo0996 <= li0996;
    lo0997 <= li0997;
    lo0998 <= li0998;
    lo0999 <= li0999;
    lo1000 <= li1000;
    lo1001 <= li1001;
    lo1002 <= li1002;
    lo1003 <= li1003;
    lo1004 <= li1004;
    lo1005 <= li1005;
    lo1006 <= li1006;
    lo1007 <= li1007;
    lo1008 <= li1008;
    lo1009 <= li1009;
    lo1010 <= li1010;
    lo1011 <= li1011;
    lo1012 <= li1012;
    lo1013 <= li1013;
    lo1014 <= li1014;
    lo1015 <= li1015;
    lo1016 <= li1016;
    lo1017 <= li1017;
    lo1018 <= li1018;
    lo1019 <= li1019;
    lo1020 <= li1020;
    lo1021 <= li1021;
    lo1022 <= li1022;
    lo1023 <= li1023;
    lo1024 <= li1024;
    lo1025 <= li1025;
    lo1026 <= li1026;
    lo1027 <= li1027;
    lo1028 <= li1028;
    lo1029 <= li1029;
    lo1030 <= li1030;
    lo1031 <= li1031;
    lo1032 <= li1032;
    lo1033 <= li1033;
    lo1034 <= li1034;
    lo1035 <= li1035;
    lo1036 <= li1036;
    lo1037 <= li1037;
    lo1038 <= li1038;
    lo1039 <= li1039;
    lo1040 <= li1040;
    lo1041 <= li1041;
    lo1042 <= li1042;
    lo1043 <= li1043;
    lo1044 <= li1044;
    lo1045 <= li1045;
    lo1046 <= li1046;
    lo1047 <= li1047;
    lo1048 <= li1048;
    lo1049 <= li1049;
    lo1050 <= li1050;
    lo1051 <= li1051;
    lo1052 <= li1052;
    lo1053 <= li1053;
    lo1054 <= li1054;
    lo1055 <= li1055;
    lo1056 <= li1056;
    lo1057 <= li1057;
    lo1058 <= li1058;
    lo1059 <= li1059;
    lo1060 <= li1060;
    lo1061 <= li1061;
    lo1062 <= li1062;
    lo1063 <= li1063;
    lo1064 <= li1064;
    lo1065 <= li1065;
    lo1066 <= li1066;
    lo1067 <= li1067;
    lo1068 <= li1068;
    lo1069 <= li1069;
    lo1070 <= li1070;
    lo1071 <= li1071;
    lo1072 <= li1072;
    lo1073 <= li1073;
    lo1074 <= li1074;
    lo1075 <= li1075;
    lo1076 <= li1076;
    lo1077 <= li1077;
    lo1078 <= li1078;
    lo1079 <= li1079;
    lo1080 <= li1080;
    lo1081 <= li1081;
    lo1082 <= li1082;
  end
  initial begin
    lo0014 <= 1'b1;
    lo0015 <= 1'b1;
    lo0016 <= 1'b1;
    lo0017 <= 1'b1;
    lo0018 <= 1'b1;
    lo0019 <= 1'b1;
    lo0020 <= 1'b1;
    lo0021 <= 1'b1;
    lo0022 <= 1'b1;
    lo0023 <= 1'b1;
    lo0024 <= 1'b0;
    lo0030 <= 1'b0;
    lo0031 <= 1'b0;
    lo0032 <= 1'b0;
    lo0033 <= 1'b0;
    lo0034 <= 1'b1;
    lo0035 <= 1'b0;
    lo0036 <= 1'b0;
    lo0037 <= 1'b0;
    lo0038 <= 1'b0;
    lo0039 <= 1'b0;
    lo0040 <= 1'b0;
    lo0045 <= 1'b0;
    lo0046 <= 1'b0;
    lo0047 <= 1'b0;
    lo0048 <= 1'b1;
    lo0049 <= 1'b0;
    lo0050 <= 1'b0;
    lo0051 <= 1'b0;
    lo0053 <= 1'b0;
    lo0054 <= 1'b0;
    lo0055 <= 1'b0;
    lo0056 <= 1'b0;
    lo0057 <= 1'b0;
    lo0058 <= 1'b0;
    lo0059 <= 1'b0;
    lo0060 <= 1'b0;
    lo0061 <= 1'b0;
    lo0062 <= 1'b0;
    lo0063 <= 1'b0;
    lo0064 <= 1'b0;
    lo0065 <= 1'b0;
    lo0066 <= 1'b0;
    lo0067 <= 1'b0;
    lo0068 <= 1'b0;
    lo0069 <= 1'b0;
    lo0070 <= 1'b0;
    lo0071 <= 1'b0;
    lo0072 <= 1'b0;
    lo0073 <= 1'b0;
    lo0074 <= 1'b0;
    lo0075 <= 1'b0;
    lo0076 <= 1'b0;
    lo0077 <= 1'b0;
    lo0078 <= 1'b0;
    lo0079 <= 1'b0;
    lo0080 <= 1'b0;
    lo0081 <= 1'b0;
    lo0082 <= 1'b0;
    lo0083 <= 1'b0;
    lo0084 <= 1'b0;
    lo0085 <= 1'b0;
    lo0086 <= 1'b0;
    lo0087 <= 1'b0;
    lo0088 <= 1'b0;
    lo0089 <= 1'b0;
    lo0090 <= 1'b0;
    lo0091 <= 1'b0;
    lo0092 <= 1'b0;
    lo0093 <= 1'b0;
    lo0094 <= 1'b0;
    lo0095 <= 1'b0;
    lo0096 <= 1'b0;
    lo0097 <= 1'b0;
    lo0098 <= 1'b0;
    lo0100 <= 1'b0;
    lo0102 <= 1'b0;
    lo0103 <= 1'b0;
    lo0104 <= 1'b0;
    lo0105 <= 1'b1;
    lo0106 <= 1'b0;
    lo0107 <= 1'b0;
    lo0108 <= 1'b0;
    lo0109 <= 1'b0;
    lo0110 <= 1'b0;
    lo0111 <= 1'b0;
    lo0112 <= 1'b1;
    lo0117 <= 1'b1;
    lo0118 <= 1'b1;
    lo0119 <= 1'b0;
    lo0120 <= 1'b0;
    lo0122 <= 1'b0;
    lo0124 <= 1'b1;
    lo0128 <= 1'b0;
    lo0131 <= 1'b0;
    lo0137 <= 1'b0;
    lo0138 <= 1'b1;
    lo0139 <= 1'b1;
    lo0140 <= 1'b1;
    lo0141 <= 1'b1;
    lo0142 <= 1'b1;
    lo0143 <= 1'b1;
    lo0144 <= 1'b1;
    lo0145 <= 1'b1;
    lo0146 <= 1'b1;
    lo0147 <= 1'b1;
    lo0148 <= 1'b1;
    lo0149 <= 1'b1;
    lo0150 <= 1'b1;
    lo0151 <= 1'b1;
    lo0152 <= 1'b1;
    lo0153 <= 1'b1;
    lo0154 <= 1'b1;
    lo0155 <= 1'b1;
    lo0156 <= 1'b1;
    lo0157 <= 1'b1;
    lo0158 <= 1'b1;
    lo0159 <= 1'b1;
    lo0160 <= 1'b1;
    lo0161 <= 1'b1;
    lo0162 <= 1'b1;
    lo0163 <= 1'b1;
    lo0164 <= 1'b1;
    lo0165 <= 1'b1;
    lo0166 <= 1'b1;
    lo0167 <= 1'b1;
    lo0168 <= 1'b1;
    lo0169 <= 1'b1;
    lo0170 <= 1'b1;
    lo0171 <= 1'b1;
    lo0172 <= 1'b1;
    lo0173 <= 1'b1;
    lo0174 <= 1'b1;
    lo0175 <= 1'b1;
    lo0176 <= 1'b1;
    lo0177 <= 1'b1;
    lo0178 <= 1'b1;
    lo0179 <= 1'b1;
    lo0180 <= 1'b1;
    lo0181 <= 1'b1;
    lo0182 <= 1'b1;
    lo0183 <= 1'b1;
    lo0184 <= 1'b1;
    lo0185 <= 1'b1;
    lo0186 <= 1'b1;
    lo0187 <= 1'b1;
    lo0188 <= 1'b1;
    lo0189 <= 1'b1;
    lo0190 <= 1'b1;
    lo0191 <= 1'b1;
    lo0192 <= 1'b1;
    lo0193 <= 1'b1;
    lo0194 <= 1'b1;
    lo0195 <= 1'b1;
    lo0196 <= 1'b1;
    lo0197 <= 1'b1;
    lo0198 <= 1'b0;
    lo0199 <= 1'b0;
    lo0200 <= 1'b0;
    lo0201 <= 1'b0;
    lo0202 <= 1'b0;
    lo0203 <= 1'b0;
    lo0204 <= 1'b0;
    lo0205 <= 1'b0;
    lo0206 <= 1'b0;
    lo0207 <= 1'b0;
    lo0208 <= 1'b0;
    lo0209 <= 1'b0;
    lo0210 <= 1'b0;
    lo0211 <= 1'b0;
    lo0212 <= 1'b0;
    lo0213 <= 1'b0;
    lo0214 <= 1'b0;
    lo0215 <= 1'b0;
    lo0216 <= 1'b0;
    lo0217 <= 1'b0;
    lo0218 <= 1'b0;
    lo0219 <= 1'b0;
    lo0220 <= 1'b0;
    lo0221 <= 1'b0;
    lo0222 <= 1'b0;
    lo0223 <= 1'b0;
    lo0224 <= 1'b0;
    lo0228 <= 1'b0;
    lo0231 <= 1'b1;
    lo0232 <= 1'b0;
    lo0236 <= 1'b1;
    lo0252 <= 1'b0;
    lo0285 <= 1'b0;
    lo0286 <= 1'b0;
    lo0287 <= 1'b0;
    lo0288 <= 1'b0;
    lo0289 <= 1'b0;
    lo0313 <= 1'b0;
    lo0314 <= 1'b0;
    lo0330 <= 1'b0;
    lo0331 <= 1'b0;
    lo0332 <= 1'b0;
    lo0340 <= 1'b1;
    lo0341 <= 1'b0;
    lo0468 <= 1'b0;
    lo0480 <= 1'b0;
    lo0567 <= 1'b0;
    lo0587 <= 1'b0;
    lo0588 <= 1'b0;
    lo0590 <= 1'b1;
    lo0591 <= 1'b0;
    lo0592 <= 1'b0;
    lo0594 <= 1'b0;
    lo0595 <= 1'b0;
    lo0596 <= 1'b0;
    lo0597 <= 1'b0;
    lo0598 <= 1'b0;
    lo0599 <= 1'b0;
    lo0600 <= 1'b0;
    lo0601 <= 1'b0;
    lo0602 <= 1'b0;
    lo0604 <= 1'b0;
    lo0605 <= 1'b0;
    lo0615 <= 1'b0;
    lo0624 <= 1'b0;
    lo0721 <= 1'b0;
    lo0731 <= 1'b0;
    lo0740 <= 1'b0;
    lo0747 <= 1'b0;
    lo0765 <= 1'b0;
    lo0769 <= 1'b0;
    lo0771 <= 1'b0;
    lo0773 <= 1'b0;
    lo0775 <= 1'b0;
    lo0778 <= 1'b1;
    lo0779 <= 1'b0;
    lo0780 <= 1'b0;
    lo0781 <= 1'b1;
    lo0782 <= 1'b0;
    lo0783 <= 1'b1;
    lo0784 <= 1'b1;
    lo0785 <= 1'b1;
    lo0786 <= 1'b0;
    lo0787 <= 1'b1;
    lo0788 <= 1'b1;
    lo0789 <= 1'b1;
    lo0790 <= 1'b1;
    lo0791 <= 1'b1;
    lo0792 <= 1'b1;
    lo0793 <= 1'b0;
    lo0794 <= 1'b0;
    lo0795 <= 1'b0;
    lo0797 <= 1'b0;
    lo0798 <= 1'b0;
    lo0799 <= 1'b0;
    lo0800 <= 1'b0;
    lo0801 <= 1'b0;
    lo0803 <= 1'b0;
    lo0804 <= 1'b0;
    lo0806 <= 1'b0;
    lo0807 <= 1'b0;
    lo0808 <= 1'b0;
    lo0809 <= 1'b0;
    lo0810 <= 1'b0;
    lo0811 <= 1'b0;
    lo0812 <= 1'b0;
    lo0813 <= 1'b0;
    lo0814 <= 1'b0;
    lo0815 <= 1'b0;
    lo0816 <= 1'b0;
    lo0818 <= 1'b0;
    lo0821 <= 1'b0;
    lo0823 <= 1'b0;
    lo0824 <= 1'b0;
    lo0829 <= 1'b0;
    lo0831 <= 1'b0;
    lo0832 <= 1'b0;
    lo0833 <= 1'b0;
    lo0835 <= 1'b0;
    lo0841 <= 1'b0;
    lo0893 <= 1'b0;
    lo0907 <= 1'b0;
    lo0945 <= 1'b0;
    lo0946 <= 1'b0;
    lo0947 <= 1'b0;
    lo0949 <= 1'b0;
    lo0950 <= 1'b0;
    lo0951 <= 1'b0;
    lo0954 <= 1'b0;
    lo0955 <= 1'b1;
    lo0957 <= 1'b0;
    lo0960 <= 1'b0;
    lo0961 <= 1'b0;
    lo0962 <= 1'b1;
    lo0963 <= 1'b0;
    lo0964 <= 1'b1;
    lo0965 <= 1'b1;
    lo0966 <= 1'b1;
    lo0967 <= 1'b0;
    lo0969 <= 1'b0;
    lo0970 <= 1'b0;
    lo0971 <= 1'b0;
    lo0972 <= 1'b0;
    lo0974 <= 1'b0;
    lo0975 <= 1'b0;
    lo0977 <= 1'b0;
    lo0978 <= 1'b0;
    lo0979 <= 1'b0;
    lo0982 <= 1'b0;
    lo0984 <= 1'b0;
    lo0993 <= 1'b0;
    lo0995 <= 1'b0;
    lo0998 <= 1'b1;
    lo1001 <= 1'b1;
    lo1008 <= 1'b1;
    lo1023 <= 1'b1;
  end
endmodule


